�y+N   x   
                       � ����                  h��0��(
�h�����(�j��0��*
�j0����*`l�����,
0l0����,�n0���0.
@n�����.@p0����0
 p�� ��0Pr0��� 2
�r�����2`t0�0�@4
�t@���4pv0�0�P6
�vP���6�x0�0��8
�x � ��8�z0�0��:
0zp�0� :�|0����<
�|�� ��<�~0�0�>
 ~�����>��0�0 	�@
0���� �@`�0�0	�B
P�����Bp�0��	�D
����00D�                ������������������DDDDDD� D�D@@@  ��O�D @��   ��D@D @��  �  @   �       ��D   �    �  O@ @  ������DD����������DODD@              � � � � � � � � �?�?�?�?�?�?����� � ��� � ��0� ����� � ���                � ��8�� 2 >������������������� �  0��   � 𪪪�J�DD����� ? � � ?�� ���������������������ꪪ������������������������    �     �  ��������������������������������������������������������������������������������������ꪪ�����������������������������������������������������������������������������DJDD���J�D��������������������������������������������������������������������������ꫪ������������ꪻ�����������������������������������������������������￻������������������������������������?���������������������������������                                                                                                                                                                                              