��N0   x   
 0                      @ � �                       h0�0�0(
@hp�@�0(0j0�@�0*
0j`�0�@*0l@�0�@,
0l��0�0,@n0�0�0.
@n`�@�0.0p0�@�00
0p`�0�@00r@�0�@2
0r �0�02@t0�0�04
@t`�@�040v0�@�06
0v`�0�@60x@�0�@8
0x��0�08@z0�0�0:
@z��@�0:0|0�@�0<
0|��0�@<0~@�0�@>
0~����0>@�0�0 	0@
P���� 0@0�0�@	0B
0� ��@B0�@�0	@D
0��00D@                  DDDDDD  DDD  DDD  ����  ��    <�8�@ ��   ��fJ  �J   (􊐊 � �� �    @ DD     DDDDD   DDDDDD   ����  ��    ���� ?���  ��������������� ������D�����   �DDDDDD  ����  ��  