��N   � `   
 0                                               h��`��(
�h����P( j�����*
�j�� ��*Pl�����,
�l�����, nP���.
�n�����.pp@����0 r���2@t�����4
�t�4@v�����6
�v�6@x�����8
�x�8@z��0:@|����<0~��P� >
`~�����>`�p�� 	�@
����p �@��`��	�B
�����@B0����	�D
�����PD �@0
�p����P2
 r�0���������������p:
 z�0���`<
�|���                $DDdDDFDUU}U��UUUU�U��UUUUU�W�UUUU_�UUUU�UUUUUuU��UUUUU_�UUUUW��UUUUUUUUUUUUUUUUUUUU����""  DDDD��������""""""""
�
�
��ꠠꪠ
� �  ��ꠠ�� � 
  
 � � � ��DDDDDddDP   @DDDDD
� �  ��ꠠ�  �������"""" ������������������""""""" UEPTAUPD D�������"""""" "  ����� """""""���������>����'򈈈�����""""""""�U��� �U�� .� ���� ""  � �P�PEE PAUT                �������"""#""�"UKP��� U��  򰈀�U�" U  ��dDfDFDDD��������""""""" ��
� 
 �� �@ DD��������  DDD������  ����

DDdDDdDDFD @ DDDDD  D D@DDDD����""  "P� ��� �U
�
�
��ꠠ�  ��  �����  ""� ������" " """"��>�>�  ? ? �������"""" ���������"""""""���IT�BR""R%R�D��HH�E!""R&%!RX����X�T%%""!"%U�Equ�R����� PP�U�  U���8�X����"("�"RR� TU  TUPP���?�?�"">%5%_UQUU��  EU  ��  UUUU��  E  ��  ��    UT""��QUTU����""  "�� �;�T�"�B�U�� ��� � ..��U��  �����  """��  ��
�     "T�����I!RbR""R�EXD��HH!R!""R&%�EXX��XX%%%""%"��P��%��_�EE� P�U� EU���8�(�X��"("h"t� TUC QTUPT���?�?�"">"=RUUU��  QU  ��  UUUU��  QT  ��  ��    UU""��EQUE����" ""  "� �;�T�""�B�U��� ���"" ..��U��  �����   ��  ��
�  """ �IT�����"R!RbR"HH�EXD��&%!R!""RXX�E�XU�%"%%%""�� PM��!%�^wuQE� T�U�  U���8��X��"("|"t"� PTU  UPP���?�W�"">"="QUUU��  UE  ��  UUUU��  TU  ��  ��    UU""��UET�����""" ""  � �;�T�""�B�U�������" ..��U��  ��   �" ��  � ��
�  """