�G��2 � �B [� �  ��J ] � � [
   �c 5 i c [�
 w  �� � � �$ [ �  ��% O � �	 [� �           � �	 [� �           �  �                       [              [' !           -  -                     1  1 [5  5           ;  ; [?  ?           E  E                     I  I [Q M           S  S [[ W                                                                                                    [�J     �  �    ��  �
�
  ��  ��    �  ��  �    � �
 � ��  �
�
  �� �    ��    �  �    ��    � �
 ��.  �     �      � �  �      �       � �     �   �  �     �    �              x [52 ��2                    ; %  Q ;  _ Q  m _  w m  � w  � �  � �  � �  � �&J)fz*�z*�z*&
z*fz*�z*�z*&z*f*)(:)h*)*:)j*),:)l*).:)n*)0:)p*)2:)r*)4:)t*)6:)v*)8:)x*)::)z*)<:)|*)>:)~*)@:)�*)B:)�*)D:)�*)FZ)�j*�j*	j*F
j*�j*�j*j*Fj*�j)�j+�j+�Z+�J+hJ+.Z+�Z+�j+(j+2Z+�Z+pJ+,
J+<
J+(
Z+zZ+�J+�j+�Z+�Z+�J+6
j+�j+xZ+�Z+�Z+�Z+0
Z+D
J+�Z+�J+�Z+4
Z+4J+hj+|Z+�Z+�J+�J+�J+�j+vZ+�j+6Z+�J+�J+pZ+�J+	j+>
J+<Z+nj+�J+�Z+j+�J+�J+,J+.
J+�J+@
j+rZ+	J+xj+�J+�j+jj+�Z+BZ+�J+�J+lJ+:j+�Z+8Z+�Z+8
J+�Z+�J+�j+vZ+*Z+*
J+|j+�J+�j+ j+tZ+zZ+jj+>J+B
j+ 	Z+�j+Dj+�J+�J+�j+�J+~J+�Z+�J+�Z+�J+�Z+�Z+�j+�Z+:
J+nJ+@Z+2
j+lJ+�J+0J+~j+J+rZ+�Z+tj+f�*��*��*&
�*f�*��*��*&�*f�*��*��*��*��*	�*F
�*��*��*�*F�*��*��*�*��*,
�*l�*��*��*,�*l�* 	�*@
�*��*��* �*@�*��*0
�*p�*��*��*0�*<
�*|�*��*��*<�*r�*��*��*2�*z�*��*��*:�*t�*��*��*��*��4
:��6
*���Ztzv��Jv�lJ),*)n:).*)p:)0*)r:)2*)t:)4*)v:)6*)x:)8*)z:):*)|:)<*)~:)>*)�Z)@j) 	�,�J+�Z+�J+�Z+.
J+:
Z+�Z+nJ+rZ+�j+�Z+�J+�j+�J+�Z+pJ+�J+zJ+|Z+8
Z+>
j+�Z+�Z+�z,�Z+�J+�Z+�z, �,6
J+�j+�J+�z,�J+�j+�Z+~J+�z,�Z+�Z+0
J+��,�j+�j+2
j+<
J+��,�Z+�Z+�J+4
Z+,
z,�J+@
�,�J+�j+�j+lz,�j+tZ+�Z+��,vZ+�j+xj+�
�z0
�p�����0�p�����rJ���2
�r�����2�r�����t*����4
�t�����4�t�����v:����6
�v�����6�v�����x�����8
�x�����8�x���������:
�z�����:�z���������<
�|�����<�|�������"
�$
����� 
�`���b����J(�j(�z(�Z($
�(d�(��(��($�(d�(�z+"
J+�j+��+bj+b�+�Z+ 
Z+�J+`�+"J+`J+ Z+�j+���� 
�`����� �`����� �`����Z"
ZbZ�Z��"ZbZ�Z�Z"jH
zJ

	���Z�J
	zL
���	j	*H

*�
*�
*
*H
*�:*�Z*�**�J*
j+�Z+Lj+�j+
	Z-��-J
Z+�J+	j-JZ+J+�z-�Z+L
J+�:
	
J

�
�

ZJ
�
�


J�J	�L
�����jLz�����L��*4
�6

��tZ�jvJ���J).z)�:)0z)�:)2z)�:)4z)�:)6z)�:)8z)�:):z)�:)<z)�Z)>�)�Z+�J+�j+�Z+�Z+vJ+6
j+�J+�j+nz,�z,>
�,8
j+pj+�J+zJ+|Z+rZ+<
J+�J+�J+�Z+~�,0
Z+4
Z+xJ+:
Z+2
Z+�j+��,tZ+��,�J+.
z,�J+�z,2
�r����J2�r���4
�t����Z4�t����*6
�v����j6�v����:8
x����J8�x���:

z����z:�z���&
(
**
:jJ��h�
�*f:&
�(f�(��(��(&�(*�(��+��+*
�+��+h�+��+j�+(�+(
�+B
Z��D
j������	�	�B�)F
�)��)��)�)F�)�*-:-*-�*-�:-D
-�:-B

-DJ-v*4
�6
�t:��n�.
Z,
jlz�Jl�(��(��(�*,�,n
,~�>
@
*�
�:��)��) �)~�,��,��,6
�v�p�0
Jp:,�J,�Z,<
J|Z��,|�,��,6

vr�2
�r
)�)�j,zz:
jz�)��)��,�f������"%" " " f�f�f�f���!�"��������"!" " " ffff�� �������"��������" " " " ff�ff@d������ �  ������ " " " jfff��h ������  fjf���  ������" jff��nf���������f���n"�"�"�"��f��� "�"�"�  ������    ����    ���             ��������        �f������  "    �n��f�f���+�"�����"���"��"��� �f���� n��̹��"� �������        �n�f� � � � �n�f� �� �    �              �nnnf������� 戈������"      ��n�f�� ���̛�� ���������"���� ;� ������        �������� " " " "��������    ��������""""����     " "    ����          ����    ""    jff��l������"�"f��������    ff���戆��!�������� " " " "fff���f������"fff���f������)��������� "����  �������� ����  �����H��"���j  �������� ���<  �������""��  �j�ԟd�X�[d��@�j�ԟd�X�[d��@�j�ԟd�X�[d��@�����,�����,��  *�.�*�.�/�""/�  D`fLf�����tf�ffffѹ�����2nnDAԙ��fnff&n&�����If�b" D&����f"�M&�jII4�)�&ff��n�I�i�����f�b�dq�C�đę���f�� HDEDDDI�n�`nff湇�������ff�f��D�������fh�hfnjf��������jff�&�.f�������Ɔ���jfG������Df����њ5����w�w��������"tDg���aa�����"�D�of"f�jd������������&TDtDtI�fff���f����������2n.tAԙ��n�`nff⹄������f���������������f��ff����������g���a�aѻ����"�tw�w�����""DD�ff�f��n�������� d�ȊH���)�!�!H��fnfnn�)�������f�j�����Y���٦��of�o����������HFhf�ffQ�)�����fff�f�f���������f����f+�)�����fbb������.+�nff�g�o�k߂"����MM�f�n�j!�����@fhfH�ff"�"���f��f�����o������"qlH�f�B�b������������f&*fn���o�a"dbff��������ofg�o��ߟ�������nffn�f����������nGFGF���������DDDD�w�����ff�f��n��������` b&b"b"��������b"ffnf�f��������fff��o����������f���f��������"c*afjjj��������fff�f�f��������fbfbffff��������&ff*jf���������������戂����DqDqff�ojgfH�������Df�(b"�f���������� N!6ff������&&f*f�f���������f�HFJ&f�����������k�m�ff����yH�a�f�f"���I����fjf�jf���������������樈����UDwDff�ojgfH��������jf��j��陚�b��j������J��k�h�j"ff�&&"*DJ�����fa�fff����������2&&"&b&􉈉������f�f�nf��������fff���f��������f"f"��f��������"*"&&fff��������                                                ~f��������������f��ffo����������g���a�aћ����"�t����w���""DD�ff�f��n�������� d�ȊH���)�!�)h��fnfnn���������f�j�����Y�������of�o����������HFHf�ffQ�)�����fff�f�f���������f����f������fbb������.+�nff�g��o߂"���MM�f�n�j!���ٙ�@f�f�fff"�"�"���f��f��陙o������"qlH�f�B�b�!����������f&*fo���o�a"d&ff��������f~g�g����������nffn�f�n��ٛ��������GFGF���������DDDD�ݟ����ff�f��n��������` b&b"b"��������f&ffnf�f��������fof���o����������f���f�ٙ�����"c"afjjj��������fff�f�f��������fjfjffff��������&ff*jfo���������������������DqDqfg�ojgfH�������Df� f"�f���������� N�6ff������&&f*f�f���������f�HFd&f�����������k�ozff�����H�a�f�b"���I����fjf�jfo���������������������UDwDfg�ojgfH��������jf��j��陚�b��k������J��k�h�j"ff�&&"*DJ�����fa�fff����������2f&"&"f����������f�f�nf��������fff���f��������fbfb��f��������"*"&"fff��������                                                �f�f������������fo�gfo����������g���a�aћ����"�t�������""DD�ff�f��n�������� d��h���)�"�"h��nfnn�!������f�jf������������g�o����������HF�f�ffQ")"����fff�f�f���������f��f�f������fbb������.+�fff�f�o�g߂"���MM�f�n�j!���ٙ�@f�f�fff!�!�!���f��濫����o�����"qlJ�f�B�b�)����������f&*fo���o�a&d�ff��������fgf�o������������f�n�f�nۙٛ�������nGFGF��������o�DDDD�������ff�f��n��������` b&"."*��������"&ffnf�f��������f�fo��o���������ff������ٙ����"c"abjjj��������fff�f�f��������fffjffff��������&ff*jf����������f���戂����DqDqfo�ojgfH�������Df�`fb�f���������� Na6ff������&&f*f�g���������f�hFf&f�����������o�o~ff�����H�a�b�b&���I����fjf�jf����������f���樈����UDwDfo�ojgfH��������jf��j������b��k�����J��k�h�b&ff�&"""DJ�����fa�fff����������2ff"fff����������f�f�nf��������fff���f��������fbfb��f��������"""""&ff��������                                                �f���f����������fg�ofg���������g���a�aѻ����"�t�������""DD�ff�f��n�������� d�ȊH���)�!�)h��fnfnn��������~f�jf������������ff�o����������HFHf�ffQ�)�����fff�f�f���������f����f������fbb������.+�f~fof�o�g߂"����MM�f�n�j!������@f�f�fff"�"�"���f��毫����kٿ����"qlH�f�B�b�!����������f&.fn���o�a"d&ff��������fg�fo����������f�n�f�n������������GFGF���������DDDD�������ff�f�fo��������` b&b"b"��������f&ffnf�f��������f~fo��o���������fff��f��������"c"afjjj��������fff�f�f��������fffjffff��������&ff*nf~����������f���戂����DqDqfg�ojgfH�������Df� f"�f���������� N�6ff������&&f*f�f���������f�HFd&f�����������k�o�j������zH�a�f�b"���I����fjf�nf~����������f���樈����UDwDfg�ojgfH��������jf��j������b��k������J��k�h�j"ff�&&"*DJ�����fa�fff����������2f&"&"f����������f�f�nf��������fff���vf��������fbfb��f��������"&"&"fff��������                                                f�fff�f������w�ff�off�o��������f���a�aѹ����"�t�������""DD��f���~n�������� d�ȊH���)�!�!H��fnfnn�)������~ffjf�ٙ���������ffg����������HFhf�ffQ�)�����fff����f����ښ���f����f+�)�����fbb������.*�f~fff�f�f߂"����MMff�n�j!�٩���@fhfH�ff"�"���f���k����j�o���"qlH�f�B�b������������f&/fjf��o�a"dbff��������f�f�fff���������ff�nff�nٙ��ٙ���f�nGFGF������o��DDDD�������ff�f�f��������` b&b"b"��������b"ffnf�f��������f}ff��o����������ff��f�晙����"c*afjjj��������fff�f�o��������fbfbffff��������&ff*off����������f�f�f������DqDqff�ojgfH�������Df�(b"�f���������� N!6ff������&&f�f�f����򙩛�f�HFJ&f�����������k�o�k暦���zH�a�f�f"���I����fjf�off����������f�f�f������UDwDff�ojgfH��������jf��k������b��k�����J��k�h�j"ff�&&"*DJ�����fa�fff����������2&&"&b&􉈉������f�f�nf��������fff���vf����ښ��f"f"��f��������"*"&&fff��������                                                fff�f�f������w�ff�fff�g��������f���a�aѻ����"�t�������""DD�ff����n�������� d��h���)�"�"h��fnfnn�!������ff�j�f��ٙ���������ffof����������HF�f�ffQ")"����fff���vf��������f��f�f������fbb��ٙ��.*�fffff�f�g߂"����MMff�n�j!������@f�f�fff!�!�!���m��f�k����k�o���!qlJ�f�B�b�)����������n&&fk���o�a&d�ff��������f�fffof���������fffnff�n���������f�nGFGF������o��DDDD�������ff�f�f���������` b&"."*��������"&ffnf�f��������fffg�og���������fff��f�f��ٚ}��"c"abjjj��������fff�f�n��������fffjffff��������&fn*kff����������f�f�戂����DqDqff�gjgfH�������Df�`fb�f���������� Na6ff������&&f�fff��������f�hFf&f��������i��j�o�j����zH�a�b�b&���I����fjn�kff����������f�f�樈����UDwDff�gjgfH��������jf��o������b��i��ꑑ�J��k�h�j"ff�&"b"DJ�����fa�fff����������2ff"fff����������f�f�nf��������fff���~f��������fbfb��f��������"""""&ff��������                                                f�nn�n ������ f����f ������ ���    f��  		�   �f�f� 	��������nf�f��������3?3?3?3? � �3?3?3?3? � � �3f3f3f3�����3f3f3f ���� f���nf�  �����`�`��Ϡϓ?�?�?�?`�`��Ϡϓ?�?�?� ff�f�f�暹��M�L?L��f�fjf�	��������    nf��    ��fff�����������  fff������������ fff����������� ��  ff��  ����    �f��  ������  �f�� �����jn��jk򙙙����1o2ff�ff�񩙩����	�	��
���������	�	��
������ �`f`fn �� �����n̦�f�f0�0�0�0��n̦�f f0�0�0� ���������� �0� � �fn�foo ������� �ff��oo ������� �f�nffn�𙟛���� �  f � � ��  � f�f� ������fnjf����f��n�j�����fjf��fnn���隚���ff���f��������jf��f�f��������jff��nf����������f��f�f���������jjf�fff��������                                                                                                @AD@ADADDDDAAA A DD@@@D  @ @A   D�f �   � @ @Dff`DDAK��&�`�� A���� ?�??@?��� ��jff��@���� �D�?D??D?����?C?C??��@� �??�?� ��o�  ��f �DD�@33ED3D3D33Do�	f3	��i�fj�f��CC�������C�C�C�COOO�CC���fjf�?�	����LN�N�MLN�M������gkggD�@����D�D�ٱ1�2q2�1pr�q�rprf�f������������������������������©�f��`�i���fo� ������D�D�D�D�D�Q����D�����`�D`�ji�������jn�oo ��������� �D�D������������� �D�����D�D��f��` ���� � fo    D���     DA   D@�	�DAn��f�D��	 �nA�f�                                                  AA@DEADDA @ADA@   @  D A�f �  D �  DADff`@DA��@F&�`�� ���� ?�???��� �D�Djff������ �@�?A?D??A����DC???C? �@��@�??�?� ��o�  ��f ��D3D3DDDD333D3@o�	fD3	��i�fj�f��C����������OCOCOC�CC���fjf�?�	����M�N�MM�LN������gkgg���@�D�@��Dٰq�2q2�qpr�1�rprf�f������������������������������©�f��`�i���fo� �D�D����������D�D�D��D����`�`�ji�������jn�oo ������@��� ������������ ���A��D�A�D�����f��` ���� � fo    ���  D      @ADA�	�@An��f���	 �nP�f�                                                 A@A AA@DADA@AA@  @ @@A   �f �   � @ @@AQff` AK��&�`�� A���� ?�???D��� ��jff��@���� ��???D?��A��D??C??�� �@�?@?�?� ��o�  ��f �D�@3A3D3A3D3A3Do�	f3	��i�fj�f��C������C���C�OOCO�C���fjf�?�	����M��M�MLN�N�M����gkgg@�D�@�D����ٰq�rpr�qq2�1�2q2f�f������������������������������©�f��`�i���fo� ������D�A��D��D��A��A�����`�@`�ji�������jn�oo ��������� �@�D������������ ��D��D��A�D���f��` ���� � fo    D���     A   DDAE�	�D An��f���	 �nA�f� 