��N   x   
 0                        @                         h �0�P(
 hp��� ( jp�@�`*
 j`��* l�����,
�l�� �@, n ����.
�n �0�P. p � ��0
�p���� 0 r�����2
 r��� 2 t �0�@4
Pt��`� 4 vp����6
�v���� 6 x�����8
 x� � 8 z0�@�P:
`z ����: |�����<
�|���� < ~� �0>
�~@�P�`> �p�� 	�@
����� �@ � � 	 B
 �����B � � 	 D
 �p�  D                    P  EO ?UOP=���UO���� �����������
������U@����UP       �?     5              D U �E���P�U������W_����O�_�����?����?���     P  P E U�T����������������������������T�P��Q�U����������������   ��� �� _����UU� ����P �����_    ��P    ��_    W�      U UPP  UPUP      PUUU  UUUP       U     UU@    UP      @ T�T�_Q @�P����_���������������������������������U  ��U�           �     �?���� ���?�� � � ���� � ��������������W���������UU  ����UU     ���_  �������U����_�U�__�_����U��_������_��___�_U�������������UUU  ��UU      ������  ��__���_���_�__���_��U_��_��_U_�����_���  U@�UP  UU�����������������U�UUU    UUU         ����  ������U�_��UU_�UU�����U�W�_��_U�_��_�����  UU�_�UU�����_�_���_�_�_�_�W� WW��_     � ��    ������U����U���UU���U�_�_��_�U�_��_����   U@�_  P UTPPUTT P@ P  PP PP U  U@U�       U            �       ������U��������UU��U_��������__��__�      �       @�U�����U�T���������P�����P������U�    �� U          �     �����P��U��U�����U���_��� _��_�� UUQQUUUUQU P          �����_    ��P          �     � P @   ���    ��@P _��     �@P       �_� T� ��U    U UPP P U@UP      E   @PTU    P     UPUPPUEQUUPPUTPUTPUQ        ���������������� 