�y+N
  � ^   
                      � ����                  h �0��(
`h��p�p(�j � ��*
Pj@����*�l � ��,
plp����,�� ��.
`n����.�p@��� 0�r����2���� 4�v ����6@x � ���P8`z � �:p| � ��<
P�0� <0~ � � >
`~����>�� �  	�@
p�p�  �@�� � 	B
@�@���B�� � 	�D
��`�p�D�np �� 0
�r� � 2
0t ��P4
@t�� � 6
0v��P8
@xp��:
0z`��|�                d`djd�����

DDDD�����jf@fff����DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD��������f�j�f��f� ������f`j��ffj    � ��  � f�ff      �       ff     ���   
���j 	������
ffj�jjf 

����� �ffj�ff     �*�   

f��       �      �???DOD�D�DO��� ����
�D�������������������������D�D�������DDG;�  qq��3p3D D

����D:C�;

��DD����DD

���#����#�#��

��������� �D�
�.� �����
� �����DKDD

���DD�D�
 ��  

DDDDDD��  

DDDDDD�TDDDDT��bbbf`@DD���	��FfDDDD������ffD�����ffdDDD���&fDDDDDGDTDDD�� 
 DDDDDD�� 
DDDDDGDTTDDDDDDDDDEDDDDDDTTDDDQDDDDDDDD0 �0 �       �      0 ��        ��*�   (��������J�*��(�⮮���⻮����.�.�
 #��"�.��*��� ��2��������/���������#������������.��� ;���������? �Q  �DD D  ���&fD
DD       �      ff��j�ff���뙩��

�0 � 0      �     0  �      �  � �*� + .(�⊮�*)���+������������*����.�#���"�
������.��2����,���/����:�������(�����.������� �⠺������
? ��� ��D�D�  ���&fD
FD      ��      �f��j�ff���뙩��

 � 0 �0   �     0         ��   , ��*� " (���:�����+��*议*�뫪���ꢺ踫��"�*�#�����������,��2/������;������(�����,/�
���.��� �㠸����
��? ��� ��D�D�  ���&�DFD  � � ��  � � �f��n�ff��⪙鹙

 0 �0 � �      0         ��    � ��� 
 (���+�(��꫸����+
��:�����⮪˪�  *����� ����,��2��������/�������*
�����<*�
���.��� ��������
��
? ��� ��D�D  ���&�D
FD    �  �  � � ff��j�ff�����

                                                                                                                                                                                                                                                                                                                                                                                                                              