��N�x        
                                                   h � � (
 h � �(0j � � *
 j ��� *0l�����,
�l����0,0n � � .
 n���0.0p � ��0
�p���00�r`�p�`2
�r�����2pt��0�P4
�t�� �`4�vp�0�P6
�v��@�06�x@�P�P8
�x ����8�z ����:
�z���P:@| � � <
 |���0<0~ � � >
 ~���0>0���� 	�@
�� �0 0@0� � 	 B
 � ��B0� � 	 D
 � �� D0                ZPZPZPZP�����������PZPZP  ������DDDD  ������DDDD@ ���������DDDD���D�DDDD�D D@D@� �     @    �𙙙�    ffUU  ������    ffUU   �	�	�    fU        @        _____DOP���������  UU          P _P____� ������    P _P    � ��________��������__C@ O�A�  ________��������              DDDD         @ @ @ @ @ @ @ @ P  P              P  P       �  UU                QP��
�P�
j  � ���������  �� ��@ @ P @P@ @ E @    UU           * SPJPZ  ���DDDDDDDD  @ D D      D@DDDDDDPZP�`Z`Z�ᬡ���
jjP Dʦ�E `
j�
�EU� ��P DDZ ����UU 
��  DD���� TDD���UDD@_____ZRj�������____�_����������       PP         ____    ����   _   ��� _____ �������     _     ���           PP @ @ P _P@ @ � ��DDD���������  DDLD� ����� DDD�Ͽ(�O���  ( �@�@� � Ё * ��� 0�0��. .    �� 
� (rr  �� � �