��N    x   
 0                      P �                         h � � (
 h � � ( j � � *
 jP� � *Pl ���`,
`l@� � ,@n � � .
 n0�0� . p � �p0
`p�� ��00r ����2
�rp����2�t ����4
Pt`��� 4v ��� 6
 v ���6�x���� 8
 x@�p��8 z � � :
 z��@� :�| ���`<
�|�� ��< ~ � � >
�~��0� >0� �  	 @
 �P�  0@ � � 	 B
 � �0 B�� � 	 D
@�0� 0D                 � ?                <       ���� ?�@�����4��30� ��D0�?���4_�� ��� ��<�������              ?��  � �P�� Q �?_�P ���   ��`  � � ��������������*�    ?? �   ���0<� ��? ? ����� �� ��?  � < � �����  � � 7� �� �     � ��     ?����` t� �   ��4� ������ �T�� �   ��        ����  ��   �P      ��        D@D       �     � ���0 �� w    Ph���    �  DD� <����� �?����  �D�D<D��<�<� �����?���?  DDDDD@  @DD    DD        @@ D             + � * 
 � � 
    ��   &ff@       �      
� ���   ff`    ���    f�            �     ,&� �DD D <        @@  D   ��  