�Y�  �~~~~~~~~~~~~00000000000000~~~~~~~~vwLMLM���~00000000000000nkmv``wMNPPPP����MN ��00000000000000 okkp{``zPPPPP�����  ����00000000000000 pkl ~~~~~~y````wPPPPP����� �����~~~~~~~GGGGGGGGGGGGGG y````PPPPP����� GGGGGGGGGGGGGG ```xPPPPP����� ��GGGGGGGGGG<=GG v`zzPPPPP����� GGGGGGGGGG;:GG ��{```wPPPPP����� �    (   (     ��v````zPPPPP����� �+++++  ````xPPPPP����� }~~~~~v```zPPPPP����� ~~~~~~~~~~~~~~~~~~~~}y```xLMPPPP����LM{``wMN (    ( MN ```z  ++++++  v````wy````xFYZFFFFFFFFFFF}y``zFF  FFFFFFFFFF �<= �JJJJJ,,++FFFFFFFFFFFFFF ,,�;: �JJJJJ ,+!FFFFFFFFFFFFFF ,!��  �JJJJJ ,+!VVVVVVVVVVVVVV },!�����JJJJJ ,+!VVVVVVVVVVVVVV �,!�����JJJJJ(,`````++VVVVVVVVVVVVVV �,,�����JJJJJ y```xVVVVVVVVVVVVVV �FFFFFGGGGG������������JJJJJ {``w              �FFFFFGGGGG ������JJJJJ v````w+++++�FFFFFGGGGG ������JJJJJ y````z+"""+�FFFFFGGGGG(+�          {````w�������JJJJJJJ�FFFFFGGGGG +�y````z�������JJJJJJJ �FFFFFGGGGG +�y````w�������JJJJJJJ �FFFFFGGGGG +�+++++y`````w�������JJJJJJJ �FFFFFGGGGG(+�+"""+y````z�������JJJJJJJ(+�FFFFFGGGGG nkkm�FFFFFFFFFFFFFFy```w�������JJJJJJJ ,�FFFFFGGGGG okkkl�FFFFFFFFFFFFFFnkm{``x�������JJJJJJJ ,�    YZ     npikl �FFFFFFFFFFFFFFkkjm``z�������JJJJJJJ ,�  jil�FFFFFFFFFFFFFFkjkk{`z�������JJJJJJJ(,�pl �DDDDDDDDDDDDDDpkkl ```w�������JJJJJJJ ��nkjmDDDDDDDDDDDDDD kl |```x�������JJJJJJJ ��nknkjkpDDDDDDDDDDDDDD |```z�������JJJJJJJ ��plpkkjlDDDDDDDDDDYZDD y```x<=������JJJJJJJ ������������������������pjl               ~~~~~~~~;:              ~}}GGMMMMI<($$
�������������%#!�������������$ � $� � &^5�@D;�F � ���������������     ��     �� ���ֵ����� �� �4O4O4O4O� �� ���������� ��            ��            �������   ������
�����������  OOO                ���     ������  ��44444�  ��������  �� ���    ������������
����������� ˜��   �� ˜��   �������   �������    � ˜��    � ����    �        ��        ������������ �����   �������       ճ��դ�       յ��դ�   ��������դ�   գ � � � ��   �        ��   գ � � � ����������������1
NOOOOOOOOMOO������OOO 4��4 OO 4 �� 4 OO 444444 OO �4  4� OO �4��4� OO ������ OO        OOO      OOMOO    OOL�A���������������            ��  �����     �   �4444��OO�   �4�����OO�   �4�����OO��  �4�����OO����������������8��   ����������   �4 �����Ȥ�   �4��  Ȥ�   �4������Ȥ�   �44444�  ��   �������   �             �             �  ���������ɤ�  �444444444��  �����ɳ��ɤ�      �� ������������������ ������ ��ը� � ղ�� � ը� � յ�� � ը� � �  ��� ը� � � � � � �� �         �� գ � � �  �� �         �� � � � � � ������������ը�����������ը����   ����������������������������������͗����������������� �� ������4�������� ������4������͘� ������4������͘��������4��������������������͘����������͗��� ��������������������.����������������������������Ҥ� � ��OOOOO   OOOOO��             ��OOOOO        �     O        �     O        �     OOOOOOO  �              ��       �����Ϥ�       �44444��       �4��  ��       �4��  �����������������A                P � d d  C O U N T R Y   F R E S H  F A M I L Y   A R M S 	 H O M E   M A D E  B A C K W O O D S   S P E L L S    C O U N T R Y   H E R B S 	 E A S Y   A L ' S    T H E   O N E   R O O M   S C H O O L  T H E   H U C K S T E R 