�Y�
 �                ��nn��nn��������33333333��������  fff  	�	�	��ff�nfff��������f�n�f�f曙�������ffffnf湹������n�@f  �@� 	  f�nfn�fn��������ffffffff��������  ffffff  ������ffff	�	�	�	�  
�
�
�  ���ffffffff���������n�n����  ` d f�  � � ���f�f���������fnf�f�n������f�f�fnff�����������n�f�滙������30303030����������  30��  ����303033  ������     f   �������������������  � ����� ������  nn��nn  ������fffffff	�������0                              �         �                 0        ��������33333333��������33333333������������������������33333333��������                                                                ffffffff��������33333333����������nn��nn��������ffffffff����������������������������  

  

��
�
��
��
���������������������������������3�3��L��L���*����*��������������������������������}��}3{37s�?����������������������������������������Z����Z���������� � � ��� / / /��� � � ��� � � ����� � � � � � � �� � � �  / / /DDDDDDDD����������������w��ww��w��߭߭߭�������������������������������������������������""�"""*(�������;��;�������������������������﨨� ��� ��
���
��0�ps030��LL��  ����������������PPPPPPPP�������������������������������������3�3��������303330�����������f�f�f������������������������ff��nn����������    3?   �����
���������    0 0   333�333?���������������000303�����������
�




����������� � ����� ����� / /���� /������������
 
 
 
 ��������    �����oo��������������**�������������������������                ��������""""""""��������" """ ��������**��**����������*"�"""""�/�..�>���������f%f&&ffX����X�����Z������_���_���Z
����_��_�V�Gd�UudU�Ie�XV�EIET�_WU]U�]]Q�WVEv�Y�[ّfQuV�ED�P �RVP`P ���n�VQQu{]SWWU���o�o_�����ֹe�������廛�������e�o�f=V�u�]��C@�a� ��� 
!?0��,�LG"B,
�@8@J�@Ģ-8 �"<��S�  h�0P0$, 0L@f`f ` ` ��� � � ff f �� 	    ff 	 	 �	�@ ` f fd� � ����        	 	    @ ` @   � �      f` Y  �� ff���o��������?3�3�  ������  ??3�3�3���������ff�f�f� ����	� �`�`f ff���  ��ff��`fff���  ���`�`� �@����� ��f���ffff����  ����߲��f"����  ������f`ff��������ff���`�`��� � ��fffoo� ����� � ff�f� ?���� = *� ?���  =��"�� o�fo� � ������������� ���������G�G�������G�G���  ���������� ;�;DND�D�DN������  DDDD����DDDD��  ������������G�G�G�G�����D�D�D�D��� ����������  ���"�"�"��������{p{p{p{p��������ZPZPZPZP������                          ��������f�o�f�ff� ����� ```````             UU����PU_U��?�UU    U   U     T U P P U T            0      ffo�  �����`����<�*�  �:    ِ  ��`f`�f������  �t�Dt7D4�  1  ��������������  ��������������� ZPZPZPZP��������ZZZZZZZZ������  UUUUUUUUZ�Z�Z�Z�UUUUUUUUZ�Z�Z�  ZPZPZPZP������        ZZ    ��    ��    ZZ      ����*��������             �            �    �       � � �+ ? <? � < �� � � � � � � �                                                                                                 ��������**��**��������������33333333��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                