�6287	 ��;|�      � D       BD   @           (DT          �    B�@            @ U�            TUUA                QU�T  P          � QU]U@T �           QUUUPU@         �TUUUT5UAU      �  �uUT�AUC�         u]UWU@U   �    �  @QuU]�@E            0EUUWUAE           ATUUUUA@       @  <uUUT PP        �  QUUT <<     @     � EUUU               QUUU@  �     �T   TUUUP        � 5U@ �UUUP          U�U@ U�UT       UEUT UuUT        ATuUU]EUUT    �     �TUUUUQUUP          E U�UUEUUP     � A@uWUQUU@         @< U]UE�U    �      < UWUuT              UTE�U@        @  ]UUUT      P UUQUT        uT  UUUUPC       UT ]UDU�@P       UUwU]T   �    A�@UQUU@��   @  AAUTUEUT �        <U@uU]UU@           @]UuUET         PUUDUQD         UUQUAC          0T UET @       =C� ]UP �   �           WTU       @ �     UU �4       @      U�T             WUPu@            @U�D�UUP          UUQ]]UUU        @ UAuATUT@         T �@ uT@ �       T uC�S�P   @ �  W@ @E@T         T ]�UQAUU@      U@U]UTUUP          PP]UUUUT       T@ ]UT T          @  �@  @    � UUA@    *         A@UQT5UU  ��       �UPUU@�             B�                P       � �      �         �                  �                                          @                 ` )   A    �  F        EQ@      U�P�     UAUQ� �    QuWTP      �AUUQ�  �   AUUEL    @UU�    3 uQp �    � TE@�     U@W    Tu@u� �   UU]]AT   �UUU     U��      UU@3    EQUP     1EDUP      AUEU @ � 4�UQ}@UP �    UATQ   �  UUUTT�   � 4EQUPD     �T] ��       ]         U@     5@]@�     UuAUP     U@T�T    SP      UU @ UEUU@T     U@@   �P T   @ �U    *@ PA     @   � @�   �      <               @         D     GT    E��P  UQL   UA    E��  �TQT �UAtT�  AUUT 1WQP    UE   4U  UQT  5EUU@   TU0  3 UT     QP@    �TU �QQ@   LL@  UEP   Q $   0QP� PU@  �0        0     D  ��WT  �G  �U � Q@@  �ME\  EU0 @U�  �U   GE@� TT\  P0    TU �A @QUW �  T   �          �D � 5� T�UD T  TPE 0T �EP  TD�P  Z   	 ��;|�      � D           �     @       �6 f@  �       �   9� � �           d dfd         @� ��	�<             f@d&@           �  ������ ��         fBf&ffd           ������<          ffffB              �����              &fff@   �  �       ����               &fbf�@          �    ����           &Bffff�           �������      �    >ff&ffn                ��  � �    @  �   l         @       �                l                 �        �     l                 �   @            � �               �           @  �  �  @    �          ��                ��@       �       ��   �    ���     ��      @;���    �� @     ��ff      fl      �����@   ���      �fff@      �l     ;�����   ��     .�fnfd      �n       ;������  ����  �  .�fffnf@   (��� .�  ������� �������   �fff�"@ "fffn .��   9������ ��������    ff��<>bfff�.���     ����=����������     &�ff?�fffff"nff�    �;��������������      &bf"fff&&b"""f@    ������������     &f&d�&"bb"""d       ���� ؈������  �   �&bf&� &""""f`     ������؈������     &fb&`02b"""""b      ���������HH�	�     bbb""fb""""�"` �  	����������� 	�      &!!""""""!"  &      ����������� �      &"   ""!" $    �  � �  �H��� �       " �  !!"� @      �  � ���  �  �   "        f@&@     �  �  �	����    "    &   &ff@(     �( ���  �����   "" �"""�  @&ff`  �` )   `        � �     d$`     @  	�     fddf    � C����     � ff@       �� �    �bf    �   ����     fffl    @  ��   @      �        @ �     @  �  ��  �     �      @�`  @     �         `    ��    9�  f�   &` 	�� � 9�   &fn�  &`   ����   ��  &fff��.f  i���� e쉙� �nfn ��&ffB̻��  bI����fn � �"f&&!��    d����f&(  	""b3��    H����bi�   �"��&d   `���H��   ""!�""&@  $H�����  	 !!   "    @�� ��  	�       f� � ��� ""0 " @    @ '   ��    $"@   	��   � fc     ��    �f` �   	�   �  �    ��     `    �  ; � �  ��@  �  �� � ff  �  ���@&f  f�!����	�f&b� ����` ��%1"!� d�Ĉ�  
"�"$ ���        @  �� �2" Fd0   8  @�  f` ��   �fp  ��  �   �  ��@  �  ��'��	� ���dfp���9��&�f���I�  "J`��" �(� !�  `��@���   � 0 	& @ � $   �  	.@ 9�0Fb� ��@��"� ((`	 ��;|�      � D          �             U @   �         �P   �  �       VT@@   �         UU!  ?�          E UUU   ?�         U@UD ���         UU �TP  �      j�@O  �   �      �eR�� �  �     � �UUD��  ?�           eEU��� ?�      �   V�T���� ��        @ Ze�����          iUD�  �   @  @    VP � �          �E@�� ?�    �    �PQ  �?�         @ VUDDf��          VeUY��[�          �U�UUVUg�         UUUUUUU��  �      UUUUUUU�         	UeUUUYU��         %UUUUUUV��     �@    Ue�UUYW��@� �     �%UReUUUg�U�          UT�UUU��E@        %UVUeV�U�T       UY��UU��U        %UVUff��U�U   @     UY�Uu��U �    @  %UVeg�DE�V   �@    	UU�U���IY  �     UVeV`DDF$        �	UU���W�Q         UUUbU? DD@       	UUUUUUW� �       UUUUUUT@@  � @  @ �VeUU�Q   �    @     UYUUUV`@   @       �UUUUY�             &VffffP          ���           DDDDDE@             	Q        � %TDDDDDT �          �U        @ � UUTDDDDD@    �      �UU � �       UUUT@DDT  @        UUU           	UUTD DDE        UUU          UVT@� DDE   @      %UeE         � � �UTP   DDD      � �eUQ            �UD  �DE@          VQ             	�U  D@            VeD   �       @ �� DD@           eUD         �U  DD         F�U@� �         ��T    O�      @��@ �     � ` )      P @  <       ?  T       UP�   � �    � ?�U@     � ��YP�   @ <��ZP @��  ? �       ?�EP�   � E@     �fUP�    � �Y�VU   �UUUU@    �UUUU`   @ oUYUUP� �  Q_�UY�`   YG�UfP  UQ�UXU`@   YD�u�U`    �!3�RU@   DD|R"U� @   �UUU@      UUUU�   �U�      BVfX      �Q�@   DDDU�     U`     D@UU� @  � @EUT     �E UT     T   @D  IV     Q U     � P U       � @�   P�F`      @�      D  U3       ��@  �@ �   T�   T 0 H� �  �%S�@@ L   �< U�� @ ��eU��  UUW�  �AUU_�  RU]$ �VU��  �T��e �UU} UUT@  @ e�	     DT@�� @Q  TD   �D� � UP� UB    %   � P@= � �0    @@ U ! B?�@  05B  C攀  �eP ��UT �TT �VTO�T  UT  V`  ��� Q@� DEP P  DP�  @  @� �    ��P�� Y��E| a��Ue  %� T   T P � B	 ��;|�      � D    �        @  � �            �          @                                       @@ �            Q              TDDDE@                       ?�DDDDDD�    �     ������      @ ?��DDDG���          ?������          ?����  @            ��            � D?�?�?�@          ��            D@<C�@     @                @ DC���D          �?��           @DD��DE  @   @   Q=�          DDG�DDD@           �=@    �  � DDC�|DDB  �       ?�@         �DDC�<DD@   @     <            TDD| DDD@�       <      �    G�DC�<DDG�        �?�� �      TDDD@DDG�@ @ �     �=�        �D|DDDDDD�        ����?�       �O�DDDDG��      ����?��        �L�G�D�G����       ����?�?���       ?���|G�G����   @    ?���?��?����        ?���G�D���� @      ���==����        @ ���G�O���      @   ���?���          ���DO���           ��������       � �������?��  �     < ����?����        �����D����j�       ��?��+��      ?��?��F�DhD|���     ���?���:>��       �����F�DhD��     C���?��	?��  �  ���G��DDDDD��      �����?��    ��DG��DDDD�D     ?������      ||DG��DDDD||D     @ ����  �   DDG��� DD@�     ?��� �        �<?�    E  �    ?����    QP  �   D�����@� @D    ��*�A!*�  @` )       �                  @P          �  @   DDD@  � �?�     ��DD��      ?���     0 �    @�?       @   @@@ ��? �     G��D@    � ��@     DDq�D@ �  QA    DD�1D@     �1    �D�GD   ��� �   �DDD��   ��<   � ?D�D�||   ������    ��O�O��    �����     ?��tO�� @   O���   @ ?��?�    �����    :3��*�?�   �F�(N���    �)�?�  �DDHO��   ����   DD�E�    3?�0�  BD��D@      ��     DD G���@� @�A 
�i@   �            A@        C�DOЀ � O��    ��  D@ @��  D�D@ <Q    D�DB  �=   LDDp 1=<   \D|� ��  �D�  �?��  �<��<� �;;/  �HJ C�??@D�D}   ?�    �  H�� D@�0    ��   @  �   � @ D  �<  O� P0B  ��   D�D  1  Dtq@  �LDG  ���  �G�?�����>� !'��DG�����@   �� �@C�|  ?� G� LD � � �� ��=4G@| �B	 ��;|�      � D                                           @          @         
�    � �         
�$    
�    @     +�
   (�           /
�    8          /
�   (�           
�h 
�
 @    �@      ����&         @  
��j��            �&�����           @  ����j�   @        ���ꩀ              ������             B������      �   � �����`    �       ������            ������    @      
j�����            
��ꫪ�  @    @    
������       �     &�������           �����릨        ��������            )��� *����       @  ��� ���`       ���� 0����       
j�� 4*��    @     *��< 4
���� �      ����< ����        ���� 2����    �  j��� <�����@      
����   <����      
����   =+����      *�����  5*���� @    �*��� p  �*ꮪj�    @ ����   @.�꺪�  �   ����     
�����   ����     
���j�   
j���    �뫪��    
����4    
�����`@   *�����    ������    &���c@   t������   �����@4  B�ꮮ�   @����� �  Ҫ��ꪀ  ����� � � 򪮪����  j�모� � 
�������@�ꪮ��� � ���ꮺ`  
������  ���������  
���ꦚ� �j������ꠀ
�ꮮ��j���ꮪ�����  
���ꮦ���j���ꮨ  ���ꪪ�����ꮪ�  
������j����������j  *������������������ ������*�����  ��j������.���������� ��������說������ꪀ �������������������� �������ꪺ���������� *�����ꫫ��몪�����   
�����������j�����    ��������j���j���      
���������� 
��     
��������   ��@    @ 
�j���   @�   � @     ���  @` ` )   �     � �    �       
       �  /�      
  #� �   
��*        *j��      � *���      �ꪀ       @�����      ���� @    j���   �   ����     ����      +����    @������    ������    
������     *k������ @  ���ꪪ�    ��jj����   �j�����  j�� :����  ���������  	�� � *���  *j�� 6
��� *��  ���� *���� *���  ��j�
����� ����������� ��������������J������ ������ꪺ�� ��꺨����� ����������� ����������� *�j����驨*���������� 
�����j��
� ������       *�   @        .     .�  � ��    ��    ��   �� �  
��    
��  .���   ����  ����  
j����  *�ꪫ� ��*ꪨ  ��*:�� ��0���B����*j����*������*���
����ꚨ*�������*�������	������耪������ 
������ @��   0      ��
� �� @ *�    ��  ��  ��� ��� �
���  &���  ���� �ʺ���L2��
�����	��*��
��*��*ꨪ��*�����&�����(*���   ��         �(  
� &�  *�!�� ������
�
�&�2�*�*�*꺨
����
��	 ��;|�      � D                    �      �   �         @ �       @  �           �                                 �f             �����            �����o�          �������9         ���o����@         ����������  �      ȏ��o��          � /��*���         � ���� ��       ꂪ�򪂫�          ����着�`     @   ���������         ���no���`@  �       ���������  � @       �fo�no��      �   ?�������          @ ���nd        ���۹���       �   ����nn`      @    ������ � @          �fffnl          �� ��//�� �        ��n�描���n���      �ۛ��/#"�����   �  ?n��f� ��fn~��     ������" ""������   �~fff興���fff��� @ ������""�+��������  >nffffo�����ffff��   ;�������""/�������   �fffffg����ffffff�  ��������"#��������   �ffffffo���ffffff�   ������������������  ��ffffffffffffffnn @ ������������������   �no�ffffffffffo��n   ������������������   ff�&ffffffffffd�ff   ��	�������������� � &f�ffffffffff@�fd   �� ���������� ��   f` fffffffff`fd   	�� ��������  	�� f` fnfnfnf` f`   ���������   	��   &f@  �f�����   fd   �  9������   ��   fd   ffnfn   �ff  ��  �����    �  @f`  fn��l     &f @ ��    ����� �  	�  f` @  �fff�  @ f   ��  � 9����@   	�   fl   >n��      &f   �   ����    �9� � &o  � f�f���  �`   	�� 	�	���� ���   f� ��fff� ` f`  �� �� ����� ��    @ff�f@ fffn f�ff �   	��� �	���� ����  @ ff@   ffn ff @  ` )                                 =�     � ���~      ?����   �?���*P      2��    >���� �   /��z��     ?����`    @ f�g��     ����@     @���y    � �����       �fgp    ����1л�  >�f�̈�n��  9ۙ� "ٙ��  �ffx���fnd����"#ٙ�� fffo��fffn ���������� ffffn�ffff ����������fnffffffff 	���������� f�fffff`6f � ������� f fnfnf d � 9���� �� dfffd  f �� ����  � `� fff@  f 	�`����  `��&ff & � d��  @�  f�nh `d  �v`�� ��  ��ff@&�`@   �� � @  @           �   ���   ?���  � 8#� �  >���   ~o� ���@   ���  �g   �C3+� C������fe�.ff@9�������.fff�ff@�������&rfffff@�����	��@f��` 	���	�&fd @ ����&f@H	���	��``f`f ��� 0              =� ��@  �� �o�  o�  ��� @ �l  zȆ�B9�r)��&fo�f`�����&&fff`		����ff A�� �$ fh `���`fBB@� � �    B  � #� �6|�@
pd`9�٘&ffd��$f`$�$&B`��