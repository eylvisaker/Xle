�,Xp�����������������������C�s��������!2C2#���� 2�� ������� ����������������� ���������������� ���!2C2A2#!  ������� ������瀀���2��1������B倀�����C�� ��B�s���3��������3����3������"�����"  ��#����3B1�����������������������������������������@0 ���"1@0 ����耀���� ������������������	��  "3B3"�   ��     ��������ꂀ�� � �� ���� ������������ � �� ���� ������������ � �� ���� �����退	    � �� ���� ���"2C2"������� �� ���� ���������  � �� ����  �����	�   ����悀�����������	!2C3"	����������"3B1������������������� 0��"3C3"����������A�����������������2��������s��#�����   �����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                r                              `	&>	��  ��	�
T  �	�
�M �`	��	�	�- �

�
�z< �
4
 ��K ��	��	�,Z �R
��i �b
.��x ��	r�	2
]� 0
r
>
�� <
x
D�� 2
 �	t �	4
v� 2
~
J�� :
�
O�� qq{?(((@?@@?@@?@(((?{qqq((/0+,.l.l.llmoA/((q  LL L  K  L L      M    L     M LA)*yw'2%%%''wxcbA$%///31(1(13///%`&(/5-t666uze/(aR K  K J K  4789:::gfvd J K  K;<=>nihJKJJKs(/������� MA(rSW�������QPL Q��L]�UMQPJWpU VVYXs(/"#NNCNN
N

						K M  MA(rS_^kNN
NN

N


						K ML  N

				MLL�Z[

N

T
T
T			MJM~N	�J��N	 �NT}|K\NT}|JBjq(/"���������K M  MA((��^�������K ML  ���������MLL�Z[���������MJM~�������J�������� ����K���JB����j����q(/���������������������������������MLMK M  MA((���������������������������������DLMK ML  ������������������������KMKMLL������������������������MKMMJM�ö������������J�Ŵ����������� ����ʸK���ʸJ���̀����JA)*yw'2%%%''wxcbA$%////%`/47��vd�������������;��h�������������������������� !HEIHEIHEIFJGA)*yw'2w'2%%%'%%''wxcbA$%////%`                 �ff�f��n���������nnnff�f���������n��f�f@������� nff     ���     &ff&ffnn��������ffof&�f&���������fj�f��n���������HȈL�LH2!!""!D��H�H��!21"!!�������H""""""""����H���"""""""����HH��"!""""!"�H�����H""12"!��H�    1"#    L�H  � !21   f���ffff����������ffffff���������fj�f��n��������nff�n�j ������� jfn     ���     &fj&�fnf���������fjfjf�f��������ff�f�fjf���������fjfnf� ������� &&f*jf�撙������f戦������""""""���hh������"""""nn�������)""""""&��*�f�f����"�)fj�f�ffj��������fjfh(�舩��"�"� jf��������"""""jf�戚����"i"''ffnf������"""""&ff&nf�f����)�")o�o"bb"b��������"""&jffj��������������)jj�j�f�b&"�&��jf��������f�f�fjff���������������"fff�d���obb""&&��������ff�ff�fb��������f��ff�""��������f�fffb!"��������ffff"""���������fjf�ff����������fjf�fff���������fjffff���������"&&&jfjj���������fjf�fff��������n��b*!f"�������bff�ff�fb��������ff��"""��������b"!"&fff��������&&f�ff�f��������f�f�ffff��������f�fff��"������HHfffb"&f&��������b"&jjfnd���������jffff�j�����"��jff�jjjf����""��f�jff�f���������jf�fffff��������fffffffo��������&�f&ff������%""nf�f�f����"�""! � 
�  �         """ ""����������   � ��   "f &  ��  � f"f"�"f ��������"&"f"&"n������� �                 �    �              �    �  
             ��������""""""""�n��nf�f���������n��fff����i ;f� f    � 	    fbbff���++�����ffffo�bf�����))�������H�""""""������ ����f �� �    j     fbbffnf�))�����fjf�f� j����	� 	��������f&&�jfjfnfd�������""""""nn�n������"�""""��H������.""""""fbbff�jj�++�����nff�h������"""""fbbff�f��++����"��������"ob&""bbjjj�j�bf�����+)�off�"o"&��������&�"&b"jb��������of&{"2"f���)�fffoof"f��������bbjffffj��������jfjfffff��������ff"fb"bf�����))�b"�ff�����������bbbfffH��))��""f�f�d�Ȉ���"�"�"f�ff""!"��������������""ffff�����jffjfjh����"!��ff�ff�"f�����������������fff��n������jj����������fj��bbf�����))�����*jf&������������"""of���H����Y�""""of���H��"a"fbfj��������&"�&��jf��������""""j&fj��������""""jffj��������ffff"&"���������f�fj�jj��������D��H�H��!2!"!!�H�����H""12"!��������fff�f"�".ff&�������a"""                               &��*ffjf��������nfff�n������"""��������f&&�f"�"�n��f�f橙�������fi�f��n��������JH�b���f���*)�ffffnf�f����)�")ffoff�ff��������nb�"������ KY!i(Hb"�&hj���i����fjf��fnn���隚���ff���f��������jf��f�f��������jff��nf��������bf��i��f:�����bff&��n���������JH�b���&���")�fff�    ����    jfff    ����    bbjfffnj��������&&f�ff����������b"&jjfnf��������b"�ff�jf��������fffb"&�f��������ff"f�"fj�����*��fff��殖��������&&�fjf�撩��������������f&��jfjfnn�������)""""��H����H�."""""�ijf�jfj��������jjjffj�j��������fjfh�f�j���"����jf��i�i����b��f�jf�f������b)�af����b���f")(�*)�(HH���hH""�b����jf�f�fi����������f��f�f���������jjf�fff���������������f&�*����fHfbf��f�����������H�Ȉ!�"�!�f�f�   ����  jj�f    ����  �jfff�f��������"ffffo�ff������)�nb,! $ ��	ffffnf f����	�	���Ȉ��!���  " " �� �� "�    "�  �  ��  �    " ffnf  ������       �  �  �      �     �jfff�f��������nff�h������"""���hh������"   f怦�� ��  "&��*�ff����"� )������� f&&�f �nfd���� �� (""nn�n������ "��������fff�f"�".ff&	�����a "�������f&&�f b nfff�n �����"��@��� ��."
�"nn����)" �" bbbfffH
�))���"&�f&ff������%"���� "  "�" "��� "��""���"��"""( ��f������"%" " " f�f�f�f���!�"��������"!" " " ffff�� �������"��������" " " " ff�ff@d������ �  ������ " " " jfff��h ������  fjf���  ������" jff��nf���������f���n"�"�"�"��f��� "�"�"�  ������    ����    ���             ��������        �f������  "    �n��f�f���+�"�����"���"��"��� �f���� n��̹��"� �������        �n�f� � � � �n�f� �� �    �              �nnnf������� 戈������"      ��n�f�� ���̛�� ���������"���� ;� ������        �������� " " " "��������    ��������""""����     " "    ����          ����    ""    jff��l������"�"f��������    ff���戆��!�������� " " " "fff���f������"fff���f������)��������� "����  �������� ����  �����H��"���j  �������� ���<  �������""��  �j�ԟd�X�[d��@�j�ԟd�X�[d��@�j�ԟd�X�[d��@�����,�����,��  *�.�*�.�/�""/�