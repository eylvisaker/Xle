��Np   x   
 0                                                h0�0�0(
0h0�0�0(�j0�0� *
0j0�� *�l0�0�0,
0l � ��, n ���0.
�n��`��.�p0�0� 0
 p@�p��0 r0� �2
 rP����2 t0�0� 4
 t ��� 4�v0�0�06
0v@�P��6x0� �08
0x0�p�8 z0�0�:
 zP����:|P�0��<
|��`��<�~ �P�0>
�~��p��> �@�  	P@
��@�� �@ �@�@	�B
������B��@�@	`D
@��� `D                """"""""��������UUUUUUUUUUUUUUUU""!" ""��������  """"�D����� " DD D��� ]" ]W]��Uu��"""P_U� ��P��"" W"���U ] """ ������P" "  "�������"       � � �   Q]UDDDDUT��""" " " ��� ����""""   ���� � """" "  ��� �  """ " ����  """   "�         �      �  ""@@����w"" @____��U�UU  " "U �� �UU" """"����� �U]UU]_]�PU���UU" ]UU]��uP��WUQQWDTDDDUU""""P_Ո���P��"""""U׈��� P��" ""P__���U����U�UU���]]U]UUU]�U��U���]U_UU__]�UUU��UU]]UU]]]]U�Uu�UUuUU]UU]_U"  "���� ����������������""  �������� ;" "�������� "  �� ������ "" ����������� �"������"  ������������""""" ������.� """ ""������ ��������.�����UUUUUU UUUUUU�.""  ���������UUUUUU!UUUUUU�U" """"�������"""""" �������"""""" ������               @              D@UUUUUUUUUUUUUU�^