���  Xb$
  :#>                          	
       gnnrs  :9:F8L                                                     9    
*          sqgns    uicjv D0/1;1J                                                   9728L  - 
# kecffdh    mchqg�021212L                                                 !Q0/1K  )  "-	,,-.) lfdcefcp   gfdcdc�/A=/6                                                ,.Q0/4      DP�w���*  kc��cehs  iefec��2K @                !                             ",,,_a6     3</��dfe~&  ue����cfn mfefffd�I                  ",.'                           FM  ,,,._<8:  F02010�ec�)  gce�.|cet  uldde��0874               -+                           C1L!,.,-_T2J   5BMH1�dd*sg����-{ffo    E��0/2A1I                                            9D0L,[UW��_`) kh ?E2�eex{��,�w��wdco    D212/1K?@                                             C22J -V�cde��* lcn  0�efcz-.}ccefcdt     EAB>@?                                               9122M[]��def�'kedh3/�ecc,wcjtkccj                                            kp            F2/11JD0����cdx~�}dce��dedz,,�j  ideo                                           mdo            D111020�����cecdcfeffcfec�,.,-)   udq                                            u            :G12/22������edccfcdcc����,-����    tv                                                         E0/011/������effdc����.,��������                                                               F12210/������cece���.-,,��������                                                               G1/11/12���/2������������������ sr                                                             H20/11/1L?=B>/������������    rgcj                                                             F000AB00J   F1��������       gdcen             rnr                                             E1/0L =21:FLG20�������   rsqg����chsrn         lccn                                             5/01;MA>@91110/�����   kcd�������ccjt          iet                                          9:  E10B2L  D11/0I       slc���������dn            t                                          F2M   ?@ H6 F/02//@     rgcc����������ecp                                                      E//:   9 ���2�/212L   kc��d������������j                                                       D22J  F2������2221J   g����������������p                                   rq                  @5BJ  D//�������02;:r���������ʙ�����cq                                  kfeh                    ?  9010������110�e�\-�[������������dt                                  ufecn                      D202������22/�cd~,,.,����ʚ�����t                                   lcccdh9:97;:9              H012���������c��`%?���dʙ���j                                     voie��0/0/1/L             E211//������R,# E���c����AL                                       rc���1122/K              H1/2/0���������.(   F��ÿ���/K                                        lfʘ��1//6 9             5B/20/12�������+   9D��������:                                        ge�����12;<2K              ?52ABB12�����*  F/����������8:9:                                   mffʘ���0112J                 @   C2/����.(  H�����������0214         �                        ref�����/001K                     E10Y�.,,
) C��������������0L       ���                      mfcf���Ɏ000B6                     D021X,-,,*  5�������������/K      �����                      vidffcd�/I@                       ?H2bX,.,-&  E����������0226        ���                        lfdfc�021M                        ?1YSPO\,SL  C2�������//>@                                    reec�1K?5K                        5/2220Y.UM  ?=�����B6@                                      ifcc�N                             510/12//N     5/2/6                                          utl@?                              ?=>@?=>@      ??@                                                                                                        