��N x        
                                                 h � � (
 h � � ( j � � *
 j � � * l � � ,
 l � � , n � � .
�n`��� . p � � 0
�p@� � 0 r ����2
`rP� ��2 t �`�P4
@t0����4 v��@�06
�v@�p��6 x ���@8
PxP� ��8 z � ��:
0z�� ��: | � � <
@|P� � < ~ � � >
 ~ � � > � �  	 @
 � �   @ � � 	 B
 � �  B � � 	 D
 � �  D                  �uuU�UUP E@Q@U U T@AP    @ @  @  =}�U�uU  UX`QVj�U�  ��P    P
   ` 	` P	� � P  X�P  `  ZZ 
�`� P (@UPUD TUU   X`Z
   �X @UQU@UTUUQ     @�       