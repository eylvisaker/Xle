�Y�  �UUUUUEEEEEEEEEEEEEEE~~~~~~~~~~~~~6666666666nkim]]]]]]]]]]]]]]]]] 









<=EEEEEEEEEEEEEE **$6666666666 kjkkmnkm<=]]]]]]]]]]]]]]]] 				qus	);: EEEEEEEEEEEEE **$6666666666 kijklkij;: ]]]]]]]]]]]]]]] 	qquqrq	)!  EEEEEEEEEEEEE **$6666666666 pjkl pkl   ]]]]]]]]]]]]]]] 	rttttu	)!DDDDDDDDDDDDDDD 6666666666666666666666  ]]]]]]]]]]]]]]]]] 	qru

	)!DDDDDDDDDDDDDDD 6666666666666666666666 ����^^^^^^^^^^^^^^^^^ 	srq				))DDDDDDDDDDDDDDD 6666666666666666666666 	s�*$^^^^^^^^^^^^^^^^^ 	qrt						DDDDDDDDDDDDDDD 6666666666666666666666 ssss�*$^^^^^^^^^^^^^^^^^ 	


									38888888887  6666666666666666666666 	ssss�*$^^^^^^^^^^^^^^^^^ 														83888888874 6666666666666666666666(	



�*,^^^^^^^^^^^^^^^^^ 				88388888744 6666666666666666666666 *     FFFFFGGGGG  	��������			88838887444 6666666666666666666666 *FFFFFGGGGG 		�>>>>���			888838744YZ 6666666666666666666666 *FFFFFGGGGG 		���>>>>�			8888874444  6666666666666666666666(FFFFFGGGGG 		�>>>��>�			88887494444      (   (            FFFFFGGGGG 		��������			88874449444 ,***,nkkm,FFFFFGGGGG 					88744444944 oikjkmLPPPPPPPPPPPPPM,!FFFFFGGGGG 					87444444494 pkpilPLPPPPPPPPPPPM� ,!FFFFFGGGGG 	U				74444444449 pjl  PPLPPPPPPPPPM�� ,!FFFFFGGGGG 	}						 (   �     @BAAAAAA  PPPLPPPPPPPM��� ,FFFFFGGGGG 	****)@@@@@@BAAAAAA ijjijPPPPLPPPPPM���� FFFFFGGGGG 		@@@@@@BAAAAAA *PPPPPPPPPLPPPM����� FFFFFGGGGG 	}																	@@@@@@BAAAAAA *PPPPPPLPM������ FFFFF<=GGG 																		@@@@@@BAAAAAA *#PPPPPPPM������� FFFFF;: GG 	U	-----------------	@@@@@@BAAAAAA *#PPPPPPM�N������           	----------------- @@@@@@BAAAAAA *#PPPPPM���N����� *----------------- @@@@@@BAAAAAA *KKKKKPPPPM�����N���� 	*$----------------- @@@@@@BAAAAAA jijijPPPM�������N��� 			U*$----------------<= @@@@@BAAAAAA 




PPM���������N�� 				*$................;: @@@@@BAAAAAA PM�����������N� 					,.................  @@@@@B<=AAAA M�������������N 						................. @@@@@@B;: AAA                 							U.................   (   (      							................. ****								                 								U																		U����										U������											~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~}				}~~~~~~~~~44568::>HMBB!,)4LLJ1���������%$!%���������, , (� %� 3� =�C�� o)� ����������������  ��          �  ��                 �������        �444444�       ��˲�� ��  ��     ��  �����������������) 
����������    �4OOO�    �4�    �4 � ���������������   �4 � ���       ��O�  �4 �б��     �ص�4�  �4��б��      �4O4O�  �4��б��     ������  �4 �б�������        �44� ��� �O4O�        ����  ��ֳ�4�              ��ֵ�O�              �������   �������������> HHHHHHHHHHHHHHHHH� �4 ��������   H� �4  ��    HH �4 ��ȵ�����  HH �4444444444�  HH ������������  H                H                H          ����  HHHHHHHH   �44� HH�D

H   �4 � HH   �4���HH   �4���HH   �4���HH   �4���HH   �4 � H    �44� H    ���� H         HH �������HH �444444HH �ʳ��� HH   ��   HHHHHH��HHH�������������  �   �  ��  �      ��  � ��   ����� �������     ��  ��     �  ר������������         ��         ����   �������������������� ������ ��ը� � ղ�� � ը� � յ�� � ը� � �  ��� ը� � � � � � �� �         �� գ � � �  �� �         �� � � � � � ������������ը�����������ը����   ����������������������������������͗����������������� �� ������4�������� ������4������͘� ������4������͘��������4��������������������͘����������͗��� ��������������������.����������������������������Ҥ� � ��OOOOO   OOOOO��             ��OOOOO        �     O        �     O        �     OOOOOOO  �              ��       �����Ϥ�       �44444��       �4��  ��       �4��  �����������������I   
               d d } d 	 Y U M   Y U M ' S 
 G I A N T   M A R T  S L E W   ' N   S L A Y  D I S C O U N T   S P E L L S  I F   I T   F L O A T S  H E A L T H   G U A R D I A N S      T H E   A C A D E M Y  D O U B L E - B U C K S 