�Y�  ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH=�����������������==���������������=Z=�������������=====Y=�����������=Z=����������==�����������=rlllllllllllllllllllllllllllllllq=��������=prlllllllllllllllllllllllllllllqp =���������=pprlllllllllllllllllllllllllllqpp =���������=ppprlllllllllllllllllllllllllqppp =���===pppMGGGGGGGNlllllllllATTTTTTT@ppp =���))ppp<MGGGGGN< llllllllSATTTTT@S pp =���)#ppp<<MGGGN<< llllllllSSATTT@SS pp =���)#ppp<<<MGN<<< llllllllSSSAT@SSS pp =���)#ppp<<<POQ<<< ooooooooSSSDBESSS pp =���������)#ppp<<POOOQ<< ooooooooSSDBBBESS pp =�������))ppp<POOOOOQ< ooooooooSDBBBBBES pp =��������===pppPOOOOOOOQ ooooooooDBBBBBBBE pp =�������=ppps         ooooooooo         pp =�������������=ppsoooooooooooooooooooooooooootpp =���������=psoooooooooooooooooooooooooooootp =��������=sooooooooooooooooooooooooooooooot =��������=                                 =���������==���������==��������==============================��������==�������================���������������������������������������������������������������������������������������������������������mnnmmmmnmm�������������������������������g�����������������������������������������������������������������g�������������������������������<		>��������������!! 	 ��������������! "
!����������������������������������                    �          ��                          ����ɗ�                          �-��ɗ�    �������������         �-�� ��    �  ��  -  ���  ����   ������       � �� -� ��� �   �  �-  o�       �-�� -�   � Ԡ���  �-��o�       �- ��-�   � � ���  �-�� 
�       �- ����   � �Ե��  �-  o��    �  -        �������   �������    ���������   �         �-�� ��                          �o�� ��                          �-   ��                    �          ����������������������������������� [ ��-�  [[[[[[[[[[[[   [[[[[[[[[[[�<[       [  [       [  																		[       [  [       [  �4[[[[[[[[[[[   [[[[[[[[[[[[              [ �������[               [ �[               [ �oooooo[               [ �





[[ �������������[ �����[[ �------------[ �oooooo[[ ���ϳ����������� 
  
 [[     ��         �������[[[[[[[[[[[[[[[[[[[[[[[[[[�\\\\\\   \\\\\\\\    \\\\\                       f\                       e\  ��������   ��������  \\  �------� ---------�  \\  �-ȳ���  -ooooooo-�  \\  �-ȵ���� -o�

�

-�   \  �-���o- ��ɳ��-�      �-ooooooo-�  ɵ��-�      �--------- �------�  \   ���������  ��������  \\                       \\\\\\\\\\\\\\\\\\\\\\\\\\�[[[[[[[[[[  [[�����������[[��������� �[[ � � � �� � [        ��� [� � � � ��� [         ��[[[[[[[[[[[[[[�O   	  
  
         � ] j r  U N I O N   F O O D S  W H I P S   &   C H A I N S  L A C Y ' S   L E A T H E R  W I C K E D   S P E L L S        S A D I E ' S   S O O T H   H O U S E    T R I C K   O R   T R E A T 