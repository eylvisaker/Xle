��N   s   
                        @                         h`�`� (
 h � � (j`���@*
0j ����*pl`�`� ,
`l����,�n`�`��.
�n�����.�p`�0��0
�p�����0`r`�@�P2
�r�����2`t��p�`4
pt����4`v`�0� 6
`v � �P6 x`�`� 8
�x0�@�08 z`�`� :
`z@� � : |P�P�P<
P|P� ��< ~ � � >
 ~`����> � �  	 @
 �p�� �@ � ���  B � � � �  D ��	�B
�	�D
�                     ��     ���    ����    ��������������뫫������ 
 ���   �������� ��� � ����U��U U���U�U���?��>�������������������� ���������������Ϫ     ?   ? ? � ���� � ����3
�UTOU�UPO�UU0�UTUUUU?UUUUUUUUUUUUUUUUUUUUUUP UUUUUPPUUUUUU  P UUUU  UPUUUU    P U�    UZZ�     UU    UUU    UUUU  UUUUU  UUU
U   UPU
U  B���
� ���@    � � ��     U UU��P�UPUU �TE�� PET  UAUUQUDUTDPDQUU  TDUD   @   DPD@P   @DPD@D@DPUUU    UU     UU      UU         �U�   wuUUUUUZU�Z�UUUZU��U             ��UUUEU�UUUU�   P U D P P       ��              ��    � � U�UUUUUU�UUUUUUU�UUUUUEEDEUUUUUU�UUUUU�UZ�UUUUZ�UUUU�UU�UUUUUUUTUUUUUTPUPU UUUUUUPPUUUUUU  
 u   ]�UWUWUUu�]�]�UU            ] WW  ] U    
�ܪ��?�p  Pq��L�LD@  5T��PPP� � � � � � � �   ����������  UU]�]UUUwUWUWUUUU�UUUUTE�UUUUQU_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTETUUUUUUU0 �   � �0  �   0 ���  �  � 0� 0      � 0<       �000� 0    0  0 �   0   �  � 