���  �&b$
  :#>                          	
                       99   9G8:r)                                                       )      gq       rDN9:F1/1��,-,*                                              ,,��     ,w��
,*     kefp     gd�2RV/0/22Z,,-[)                                         �� ,�� �#  }ed�,,   md��hq  rdd�0YO����1W-[]1W                     ,)           ��	,,.��
�� �򍖍%     ul���hsifdcc��fec�_`,T/0Y,,,.,T8:                9,[]J93;78#      ����,������
�/�>=}n       ld���fnkfefcedfe�-,,.,U1Z-,,,.S10:              32Y,S021/0//6         "�,�����,T/�en mcdh       ie��fhldd�dz�c�Y\O^]\T2R�O^\\,V2/;8         9D//PO/0Ra/10I99:       -.[����,[�/�hskejt      kf��dtk��Y�-,�a2/112YT2^]21/Y.U//11X#      ���0//0/ZU0201YV28# #  UR,[\.U�/�ecdj        le��j ?0=2^SP-O22221YS0/211//P1101/P�      ��Q//1/6 G/1/01ZV1/K # ( CR,[X,Q풓ef�o          i��n  ?=A5/P]02/22/02/12210/01/00/��-'     ��._a/>@ G�2/02Z_0I  ) "( CW,UX,Q�ede�$��        ut  gcnF012101/2202/11110020/�/1��-+   .��,    C�10/R`O0J      !`OZ-,}ec�������            mfdo F20100011/110/2/0/0/2012/W-,(   ".-��      C/00R-,1024      ��,ZX,|fd�//�����      34: kej sC222///0/11//0RT10222��1��    ,,��     �!V1/P\,V/Zb97��S0^\O��00�����       ?H1K ut l��1//R_Ta/0Z`QR-U0/ba0/�1��      O1��    ���O1�/2P_b`.,���U���O/b[//101����     #  @       mce�02X,,-Q1X,,-,22b`,_Q//6      !221��   �������00/W,,,,�������/2XV022/20��      9   �rhsrgzzQ/b+aX.,,-QZ.-,��1K    -Q22��:�������Q/�`,.-,����2//��^U01001���      !.,T88�����d���-%@   ��W-,,,,,.�����@ F87\,OWS//���O/L  "��,���������-,V0/�ef�0/RV/�cfo     .,-T0�����,�,,,,,)  � ���Y�,.,,,�����   E1/WS1XS1���022@  ���,���������,,T/�fec�0/P_0�cen      �,[Z��������,.,+  ����������.,������   G/2YU2YU0���/2I   ��,.������,{���wdcd��V00bS2�fj  9     .TX��� ����(  �����?����,����&�    51=01ZQ�2�2��R
)���,,������,|dffc���,SXV1PO0At  3/4 8# ����   �        ���  ���,-����  ��  ? 21X,��/22��,)���,,������.,,�cc�,.-,UY_a1/0K  F11M!S/8# "�����  ��        EJ ����"����� ������QR.����a11W,*����������.,,-{dc��,,T�R,.V/1L  D01J"U16�:!������ ��       ���������������� �������������S2/Y,,����������-,,,.������}c��._V0J  5>@@E1RQR.-�,,����       ������������������   �����������211P,,,���������.,-,,,,����cdd��_02L     FZ.,�-��-,����������������������������������������������.�����������,,,�������efcd�S/I  FL   5W�������������������������������,���������������������������,�������,��������d�ccU2�� DJ    "������������������������� ��������������������������-,�����.,%�     �������������Q��� C24  !���,�������.�������������	������������������������,,.,������&     m�ʗ�����������,V�� 5/1K .,,����,,,�,,-,,����,,-���������������,����������������,,,,-����'      uiʗ����������,T6   H/4,.,-����.,,,,,,,.,-,,,,����������������-�������,,-,,,,-.,,,.,,,-,       uʚ�ʗ������-UL   5/I ���.,,,,,,,,,,,,,,.-���������������,-����,,,,,,,,,,,,,,,,,,,,.#     kc�dc������-S/4   92K �,��,,,,,,.,,,,,-,,-,,,,,,,���������,.,,,,,.�,,,,,-,,-SP-,,,,,-,)      vide�����.�T1J7L9D0J.,,���,.,-,,,,,,,-,,,,,,,,,,-,�����,��,-,,,,,,,,-,,.,,,-,S0P-.,,,,,'       kddʚ�~-.,T11/12/2I�,���,�,,,.,,,,,,,,.,,,.,������ႂ�.-,,-,,,,,,,,,,[]\,\U2/Y,-,,,       lce��c���O001/001M!�-�"�����,.,,,,,,,,,-,-&�}ffex��}fd�,,,,,,-,,,,,,,,S/^O00/01P,,.,)��       lcjutv�����//��/A6,,�,,.�,,,,,,,.,,,,.,,(kddfddfffdfddx,.,,,,,.-,,,-U//0////00/X,,,
���       v     �� D�����   -".,,,,,,,,,,#geecefdeedccde�w�~,,,,.,,,]2001//0//1����.,���             ��F/����        �    ,mdedcceedefdecefcd,,,,,,,U010/20/1�/��������,)            �?@��          ���      ",(      lcfeeeefdfeddffec�,,,,.,,T///0/000/��///�����Y]L                         ��  ����� �  !$#   rq g���fdededeeefddz,-,.,,,,,Q012/00/0���20�����/R'  �                     ��  �������     gffd�����fdccefedeed��,,,,,.,,S000/000����00/����0Y.,���#  )                ,�,,,(�     ude������cfcefecdeffff���.-,,.S00//0/0���00/00//0/Z,,������,-(          FK ,,���,$�������;��������eeecfcffddefdfedx�}~,T001/�������1�2������,�,���& ",.,* *        F4����,��������/R�������e��ceccfeddtuiedcfdo-Qb`�����������������������	,.,,-	�#        D/L  �����,.������b`,,-,-.������fcceffep kcdffj  .,.,,-�������������/���������,-,.,,.,       G/8: �������1Y\[]W.,,,,.,�������deedech ljvut  ,-,,.,������������񑋎/�����Y^\-,,-,,.-)      ?=R`-)������/1/00b`-,,,,,,��/A����e�ddfden       ,,,,�,���,-��/1�fc�/11��011Y,,,,,,,,*        -,
,�����/2/10Y-,,.,,,.T/N H�����efecj           -.,,-.�,,���00edd2/2//012/2P-.\-,,%        ",,,.,�����//220\,[\,SP\��1KC����cceco            ,*"����,,-��cc�101���10021WS2P,,,        ,-,,�����0�b//Y.SPO20/��/M����fdfjt #           ")��.,,,Q�ddcf�10����02100YU0Z,-         ��������X����,TA@=/2//0/���cccn   -(               �,,,-.}ec��ed�0����/11/0//b`,-)           ��"���������--   G122/2���dceo 	-)            ,-,|fd�1/�dc���0/2/1X`_`,,-,.*            ��������� 977/1//1//2�ddch� .,*         -,'  ,,-��0202��0�100011P]W,..,-,&         #  �  �� "��(9<;2/00///10��cc������-        �.,#  ".,,,,V1����/0�0/1110122^\\.,,'          #   ��  F02221/1/21210�c�.,����+          ,-    ,.,,.T10��/2//0/102/02/20W--,-(         #) ,)     ��200020///1/�fd�����           -,,,,S�����1/10/101002ZT1Y.-,,)        @ !-
	.
����00/02110/21����������             ,,',,,-,������Q0Ra10011bVXO1Z..,+            ,,,.,,-,���,�2///20020/11222�� ����       ,�#  ,.& .,.,������,`-,/2110X-_00X-.,(            -��.��������0b21200//2/Z`����� ����������.,) �!.,*,,,-(������_`,O///0R[^]/ZX,,&          ,��,��������@V201201//P,,���� �����������,,*���.,-)  ��,,[PO1/110YU2/0/]P(         !,,.-���,,�����    �/11/1010Y.�����  � �������,,����,,,*        ".-T///22/1/1/0/11Z*          ,.,����������������1/120111PO����������������������,,&        _a/1/1/22/2/000Z.     ,�������,,���������///00120222�������������,���������*           "._Q0021111/0/b`-,,,'        �������,��1022/��01100122100/02Z.,��������,�,,�����'           ,.T012/20211R.-.,,.,'    F874 ������,.����/����T0112/1/22122���}~������,���������$ss       !-[]0/01///1R.[\,,    D0`:����������0����U2002/011/20�dcedd���,.�����������{���dh      ,,S002/0210/Y\O1^O4:      F/0P,,U/���������20/���210210021120�eeededdd~.����,������|d�|cdn    --U0/00/0/1//000//0J     ��22PO/1�0��������������211//012/1R|dfefez��,,,����������}f}cehqkqrgx�VRTRV01001//1//Za6     ����11�������������������010110/0b`,weecfd��,-,,,,,��,,,-{�f��ecd����c�������/0/01����/R-     ����2�����������������/20122110X-{ceccfc��.,,-,.,,,,,-,{f����ce������������00/0�edc_-,,,)   ��,_Q�����������������10��2���/Y\|fcc���,,,,,,.,,,,,,,|������������������U/����cc�/W[]/P(  ����,,,�����W,,[\V0�-���_a2�e��fd�22W�cz,.,,,,,,,,,,,,,,,,,������������������U/�efd��10PO10Z  ��.,,,.,�����,.TY,/W,,,,-T/0fdced�/1Y,,,,-,,,,,�-,,.,,,,�-.������������������0/�edd000///0/X,) ,,,,,,,,�Q�X.,UYO2P,,,,[]02�d������X,,,,,.���}d~,.,,,,��,�����������������ʣQ��cd�100/��/0X.*  ",,,,,,-,,�,,,Q11/R,S\,T����fe��cce��,,,w�fc���Y\-,.,,��.�����.����������cc�}dddc�1//�������,( 	,,-,,,,,,,,,.S00Z,-UX.T2�eddecdddfc�.,}ecd�0121XO^OW,,,,.-,��,����������dfdcddcc�//00/0����� ,,,,,-,,,,,,Sbb`,,_`,[b`y���fffecfx,|fe��/0212Y22/X,-,,��-��-����������dddeeffe���110/Y-��    -,,.,,,,,,,,,_,,,,,,,-,���U1�ec��edc��|�Q022//020/0^^\,,��,��������������e�|dcecdfd�//���'��  ",-,,.,,.SW,,,,-,,-,,,.{fdd�1�fe~|fdz��,,S/12220/12/01W,-.,-���������������,yecdcefde����� !	,.,,,[]2^\,,,,,,.,,,|ccf��dfd�}cf,,[]/021/0220101/Y,,,,,��2��/����������,.�dfcdcf������'  "+ �-,[]0102X,,,,,,,,,,,�fffcz�����f�~.T0100RQ010Za/02Z,,,,,��/bQ2����������,.|���yc�����    ( ,H2//1b`,-,,.,.,,-.,�df�-.,,S�cd,S121Z-.a2/X,V0R.,,,-,U/X,,V���������,-,.,,-,�,���(          U20/0Z,,,.,,,,,,.,,-��\,,,-]/��,,O22Z`,[\Qb`,_aPX.-,,\OZ,[]0Z�������.,�.,,,,.-,�����       =22b``,,,,,,[]Y,-,,,,O0W[]]0/2W[]0//X.,U0P\,,,-.,,,,S0b`,T01^\.,,-,,-,,,,,-������������)      F00X,.,,-,,.S11X.,-[O12XS0/2/020/2//X,T2/2X.,,.,.--,_b`,,,U20Z,-,,.-�,,,,,,�������������   *97/R.,,,,,,,,T22Y,,[0/22YU/N?@=A@H10Z,-&C1/X,,,,,,,,,,,,,,,V22W-,we�,-,,,�������������   ,,TR`,,,,,,,,,,S0/R.,T//N@5A?@     !V2X,.*EA6,,,,.,,,,,,,,.,_a/Y,&  mddf��'��������}�q   !,,.,,-,.,,,.,,-T10X,-.Q1J          Tb,-,'   ,,,,,.-,,,,,,-.,,,.-(   vicep  ��,������dt97<X,-.`,,,,,,,,,,,U01P^[UJ          "-,)  !,-,,,,,,,,.,,.,,[OZ,)     uehq�������쒓~}dnD02Y\,,,,-,,,,.,,.O121/2^K ?@              (  ,,,,,-,,,,,,,,,[]/0X,*     gfc����������cejo D/2R-,-,,,,.-.,,,O21/20/2K                      -,,.-,,.,,,,,-.T22Z,-&     tf�J    �  ��cco  5/1YU^-,,,,,-S0/20>B06                       ,,,,,,,,"&U012^\*     m�A�   rq  ��dj    H2/22J ",,.,-.U/2N@  @                           ",,, 5/0//Y     @  rqkceh ��uv     F22002K -,,,?=>K                                   ,,-(    @C01N          idfdfcp          C>B6@                                           +       5>@           ljutv          (%@L+%@#KU+5JW5N 0L )DP8Z*"<]ZRIPbb BN CPN>@>	>	1?5&L 0 I8	W]DZPNQ	0>H:B 6& cU4>^ ::F_\	?  AQ:F,0b	P90Q! 2K _V 	G6V;1A^@FQ-/ JF QJ.>]	!Z%!]'% ^` %E=JB.DXb	I3-:>  5F5F]4KV4Y0 > >0_UZ%UZ%MPRZT +V 7 	WRZ)_V_V	:="W0I:; (1 CPZR	R	P@`/=@ > @#_0(7?2,:,:X
 K NQ NQL.<@TKW38#@B8# ? WbcK) ) IUIUIU ^ %<	C<	CEUE-b4b4"T ?0 ]]:;P?(PE' $] $][H"D][H"	 6'" =I []?0/[]:[]:]:',"," 5H #5H\5H\)I#@OOK L FWFW22.\MHH2Z 	 	T'2[>1_	c2=I_?=I $ B_	TDYDY2`D22 = =