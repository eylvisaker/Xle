���"+�7                : :: :    ::::::::::     : :   ::::::::::    : :  1  ::::::::::  1 1  ::   0 ::::::::::     :: ::::::m::m::8988988998989888 ((8) 9)*8 *9++ (89)98  (  ).)88(.8998*89+*  +  99/+98*/*85959(8 * 5 5 ((9,8,9*88+94949)+ 4 4 ) 8)9-8-9+:;;8<:8<=9:=8>>::?:;:=:?:8;9=9:8@:<:>:@:8:9<9>8::::;::<::;98<:89:=::>:::98:=89>:ABBAAABBBAAABBAB $$B% A%&B &B''  3 $ & 3 3 32 % ' 2 2 2   %  $  '  &    :CCBD:BDEA:EBFF::G:C:E:G:GCBH:D:F:H:AFH:::DJ::JCD:BCFI::IE::IB:E8KKBL8BLMB8MBNN88P8K8M8PMB8PO8L8N8O8O8BL88LR88RK8KRBNQ88QM88BQN8STTSTTSSSTTSTSTT:UUSV:SVWS:WSXX::]:U:W:]:]US^:V:X:^:TX^:::V_::_UV:T_X`::`W::`T:W8YYSZ8SZ[S8[S\\88a8Y8[8a8aYSb8Z8\8b8T\b889Zc88cYZ8Tc\d88d[88dT8[BeeSfBSfgSBgShhBBiBeBgBiBieSjBfBhBjBThjBBBfkBBkefBTkhlBBlgBBlTBgnnonoonnononnoon   n! n!"n "n##  7   " 7 7 n6 ! # 6 o#6   !   ! o#  "  o ":uuoo:oooo:oott::qno::nqonp:pn::nro:r:o::oso:n:s8nonn9onon9oono98vvnw8nwxn8xnyy8z{|}~����������������������������������������������                             �               �               �               �               �               �               �                          0               0               0               0               �               0               0              P      UUUU      P      �* �    ��            
(    ���      �     PZ�     
Z      ��	�    ff            ��    `df UUU UUUU@ P U@UUP T UTUUUUUU UU U UUU@U U UPU U@P U U U UU  UUU@U@P U UPT T UP  UUUUUUPUUUUUUUUUUUUPUUUUUU     UV  QUUV  T U@TPP E UP�TYUQ U U  �UU D � QPT T      
��  �
��  � � 
�  � ���*�*

� � � "  *����   � ���      � � �  ff  �  � ` f f`f`	� � 	f f f  ����� � f`f f   		 � ��f f df��� � ��f f F f`  	���� ffdffF������ 	dfFff  P U U P U U U P   U U   U  � � � � � 
�( �   * � 
 
 � " �  � � f F f `  	  �   f f  � E Y P U U  P   Q �  U U T �������FfdfdfFf������dfFffdFfUUUUUUUUUUUUUUUUUUUY�U�UVUfVfVFUU�U�U�eUfUFefeY�Y�U�UYVfUfUFUU����U�UfefefUUUUUUU�UUUVUfUVUUUU�UU�UEUfUfUUU*����
��

�(��*�����*�


���UUU�U�P�UZU�Z
�
UU
U
U��U�U�����
Z
U
U
`�U�U`UU���U���U�
	UUUUZU�U�U�UZU�U
UZU�U
U��%U�U�U�U�*R�UUUU��jUUUUUUUUUUU��UUUUZ��
�� ����f*`�j
�
���������F
&
��
��������*
F�f*f
����()��*
�f���f!��*���f�&�d�F�
�����fbf(j*fb��� ����Hffdf������Ffff&������������������������������U]U_W���U�U�����UU�U�}���U�U������W�WU__�_�U^UW������U���U�UUU���������of�����ٙ�����n����������������g�f��������������nfU_UW�WU_U�U�U_�U�U���U�U�����UUUUUWU_�UUUUU�����u�UUUU��UUUUUU���������o���f���������f�f�f�F���������f�f�������������ffoff慠�.���㨠
?�����������
���
�*��?������

������������*�
�
���������
�
��
���������
���
�
������着

������������
�

�
UuUUUUWUUUuUUUUUEQYUQTUTUYTeQUUTeVEUEUTEUU�UE�UUUUUVUEUUUUUUUUUUeUUUUUTUUEUEU�UUUTUQUUUUTUQUUUVUUUUEUUTEUEUUUETUVUUUUPU�UTUQUUUUYU��E�QUfTeTfYUQU�XIUYUQFfVE�TU��U�UY�etfEffUUYU�E�Y�E&TfFfEUUUUU�UUUUZU�U�UUUU����UUUU��7�U�Z���U���p������_�_�Z��_�UUUUUUUU@UUUUUUNUUUUUUUUUUUU��K�@�TT�N�T�T�T �������. UUUUUUU�UUUUUUZ�UUUUUU�UUUUUUU��������UU������UU����UU���UU

���� ���

�
��

����
���

������������������
���������EVQDUP  UUe@ �UQU  U��   �0 0ET   UTU   VE�  �UQUUUUUU_U�UUUUUU�UUUU_U��UUUU_���U�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (                        P  TP  @  E   T@   T QU EUE  QU  �  U   U@  AP   P   T                          (  �������������������  ��  ��� ��� ?��� ��   ��   ?�   ?�   ��  ��� ��� ��� ���<�� < �����                    (                        �   (   �    �   �   ��  "��  ��(  ��   �   ��  ��  ��  �(  * �                          (  ������������������������� ���� �������� ?��� ��  ��   ��   �� 3��� ��� ������ �� <�����                    (                  p      p    �   t7@ ��� G4 �  44t4    w              ��                          (  �������������������� �������  ?��  ��  ��   �    �    ��  0��   ?�� 0��� ?��� ?��� ?��� ��� ?�                    (             �      �   ��� �� ��� ?����?���0����
������ � ( �  ��  2��  <��  �(� �
?                          (  ������� ���� ?��� ?��  ��  ��   ��   ?            �   �  �  �  ��  ��  ��   �� � ?����                    (                             �    �    �   �  *��  ⨯ Ĩ<  �   �   �   �  �  < �  � �                          (  �������������������������� ���� ��������  ?�   ?�   ?�  ��  ���  ���� ?���0���0�� ��� � ����                    (                   0      �� <�  8   ..   �   ,�  �;8   .,   �         �    	�   �    �                         (  ��������?�������� ���?�?���� �?� �?��  ?��� ��  ��  ��  ���� ���� ���� ?��� ������������                    (         �(   ( �� ?��� ��� ��  ��������?���0?( ?�� �� �<� ��?  0� �� 
< ? (�?�                         (  ������� ��  ��  �   �   ?�   ?�   �               ��  ��   ��  ?� �?� ��� ? ? � ��?�?                                                                                                                                                            � � !�!�!z"?%�%7&�&/'�''(�()�)*�*+�+,�,�,{-�-s.�.k/�/c0�0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (         w   ��  ww ]U  wT@ ]P  u  ]D  uE@  ]@   WP   P   T    U    PP   U@    P                              (  ��� ���  ?��  ��   ?�   �   �  ?��  ���  ?��  ��  ?�� ��� ���� ���� ��  ��� ��� ���������                    (           @  P@  @  p  �  Cw  ?�  �0  ??�  ���  ��   ��   ?�   �   �    �    <                          (  ������?���  ?�   ��� ����?�  ���  ?�   ��� ��   ��  ��0 ��� ���  ?��� ?��� ���� ?��� ������                    (        	��  `     �` `� � dfb@ ��� ddf  �  $bd  ��  Fd  	��  &f  ���  Df@  	��                             (  �� ��   ��   �   �   �   �   �   �   ?�   ?�   ��   ���  ���  ?��  ?��  ��  ��  ��� ����                    (          0?   �?   �3� �3� �<� <<� <3< �3? <�<��3<���<3��0?�0���� � <0 ��� ��                          (  ��������� ?��  ?��  ��  ��  ��  ��   ��   ?           �    �    �    �    �   �   �   ��<?�                    (              " �"" ������  �(( 
�      �   �� 
��      (  
�   � �                                    (  ������������������?����? �  ? �  � � � ��   ��  ��  �      ?   ��  �� <���?����������������                    (          �   (   �    
    �(  ((���
((��
��*�" ���("�� *����
��*  *���
���� *� �
                                 (  ����������� ?��� ��� ���  ��  ��  �    �                �   ?�   �       �  ��?�������                    (            < <  ��  <<       <� � �0 �  �;�  ?�  ��  ��   �   ?�   ?�� �?���?�                              (  ����������   ��� ��   ������ ���?�� ��   ?�   ��� ��� ���  ���  ?�  �  �   ?��������                    (                  � �  �   < �   p � � t p ��� 7t  ��@  �pt   4    � 3@4 � �  0                            (  �����������?���� ��� ?� ����?�����  <�   �   ?�   ��   ��   ?    ?    ?    � ����������                    (       0��  ?*:� ?*�  ʪ�  �  <*  
� *� � * �� *��� 
�    �   ���  ��� ��  � �    � � *                          (   ��   ?�   �   �   �0  ?�0  ?�   �   �   �   �   ?��  ?��  ��  �� 0�� ���� ��� ?�?���                    (               8   � �;   � � ��,�� ;�� �.�  ���  ..�  ;��� � � � � , � �    ;�                          (  ������������� ����� ?� � ��   �  ?    ��   ��   ?�   ?�   �   ��� �0� � ?��0�� ����?�                    (                  �    �   
��   �   �  ��  � (   �   "    �  �   �         �                                    (  �����������������  ��� ��� ?��� <��   ?� �� ���� ?��� ������������ ���?�����������                    (        �    ��  <��  �� ��� ��� ��?����?���?0� �?<��< ? << ��<<��< <<��<����    �                         (  ��?����?��� ��  ��   ��   ?�   ?�   �   �                           �    �    �   � <����?                    (         
�  ��� *�*� ���� ������ʀ�*( �*�  ���� ��*� *���  ���   (�  ��  ��� *�� ��� 
�                            (  ������  ?��  �   �   �   �   �   ?�   ?�   �   �   ��  ��  ��  ��  �   ?�   ��  ��?���                    (       �  00�0 0� �  ?�  ���/0?����/ ���  �� ���0<�0�3�  ��  ��  ��  ?��                          (  �?�����?� ���� ��  ?��  3��  ��   �   �   ?�  �<0  ?�      �   �<  ��� ��� ��   ��� �                    (             *�� ��� ��� 
(�* * �  ���   �� ��� 
(*  (   � � �     � �    �    �                         (  ������� ?��  ��   ��   ?�   ?�   ��  ��  ��   ��   ? ��?����<�������?�?�����?� ����                    (                       �  ��?�  ��� ���0����  ��0 ��������Ã�< ��  ;�   <0  �   � �                              (  ������������������?��   ?�   �   �   �   �   �       �    �<  �� ?��  ������ ���������                    (        � < ��  � ?  ?��  ��   ?�    �  3�   �� �   <0   � �   ��  �   < <   �   ?�  ��                         (  �����   ��   ?�   ?�   ��� ���  ?��  ��  ��  ��  ��  ��   �� ��� �� < �������  ��� ���?                    (                   
     � 
 �(  ��   "    ��  ff  	��  ef@ ���  ef`  ����ffd  ��� `    �                          (  ������������������?��� ��< � ��� ���  ���  ?��  ?��  �   �    ?�   �   �   ��0  ���� ?��� �                    (             T   HQ@  %P  �T  T  PP   T       A     T   P   QP  @  @  A                          (  ����������  ?��  ��  ���  ��   ��� ���  ���  ?�   ?�   ?�   ?��  ��� ��� ?��  ��  ��  ?��� �                    (               �  
�  (( �H@ 
!!  DDD@ DD@ B�D(�  D�! (   DB    �    �                              (  ���������?���<��� �0  ��   ��   ?    ?�   ?�   ��  ��  �   ��   ��   ���  ������������?�����                    (        �   <   0��  (
   
�<  ��  2�  ��� ��< �?? 3�< ?�� ?��� ��� #�  ��  � � *����                         (  ������ ���  ?��  ��  ���  ���  ?�   ?�   ?�   ?�   ?�   �    ?    ?�   ?�   ��   ��   ?    �   ?                    (          0        <    �   �     ��    �        <    �   � �?� ��� <���0?�<0<��000�00                         (  ���������������� ����������� ?��� ��� ���� ?��� ������?���  ��        �       ��?��                    (        �   8�� "��. ;������������ �  �  �  � �;�������;����.���;� �,   ;  8                          (  �� ���� ��   �            �   �   �   �   �   �   �   �             � ��? ?� ������                    (       ��  <��  �� ��0�< � � ?�������=�����<�?|<�<��<�  < �  ��  � � <  0  ��                          (  � ���  ?�    ��   ?�      �  �   �   �    0   � � � 0? � ��� �� < �� ? ��0? ��� ?��? �                    (        <   <��  ��  <�   ��� ��� /�;�   <��  ,�? ��� �Ͽ�?�� ;�� <��?��� � ��� ,   �                          (  ������� ?��  ��� ��  ��  ��   �    ?�   ��      �   �   ��  � �  � �� �� ?�?������                    