�7�  (0
�
0�p
�
p�    0�0�p�p�    0�0�p�p�    0�0�p�p�    0�0	�	p�p	�	    0�0�p�p�    F @ �� �     @     r�
�                                                                                                                                                                                                                                                                                                                                   �((�                                                                                                  �  ?�  �� �� ��  �  ?�  <�  ��  �< �?     ������?���?��������  ��  ��  ��  �� �� ��  ��  �� �� ?�?��              �  ?�  ��  ��  ��  �  ?�  <�  <?  � <     ������?���?��������  ��  ?�  ?�  ?�  ?�  ��  ��  ?���� �?����              ?�  ��  ��  ��  ?�  �  ?   ��  ?�  �  ?      ������?���?����� ��  ��  ��  �� ����� ?�� �� ����� ?�����              �  �� ������<?�� ?�� �� �� �<  <   <     ������?���?�����  ��  ?�  �     �  � � �� ��? ��� �����     
         
�  :�  �� �� ��  
�  *�  (�  ��  �( �*     ������?���?��������  ��  ��  ��  �� �� ��  ��  �� �� ?�?��     
         
�  :�  ��  ��  ��  
�  *�  (�  (*  � (     ������?���?��������  ��  ?�  ?�  ?�  ?�  ��  ��  ?���� �?����     
         *�  ��  ��  ��  ?�  
�  *   ��  *�  
�  *      ������?���?����� ��  ��  ��  �� ����� ?�� �� ����� ?�����     
         
�  �� ���
���8?� *�� �� �� �( 
 (   (     ������?���?�����  ��  ?�  �     �  � � �� ��? ��� �����      �   �   �  �  ?�  ?�  ?�� ?�� �  �  ?<  ?  <  ��    ����������������  ��  ?�  �  �� ?�� ��  ��  ?� �?� ���?      �   �   �  �  ?�  ��  ��  ��  ��  �  ?<  �< �0  �<     ����������������  ��  ?�  ?�  ?�  ��  ��  ��  ���� ��?��      �   �   �  �  ?�  ?�  ?�  �  �   �  �  �  �   �     �������������� ��  ?�  ?�  ?�� ������ ��� ?�� ������ ����      �   �   �  �  �� ��������<�  ?  � <� < � <      �������������  ��  ?�  �  �   �  ��� ?�� � �� �� �����      �   �   �  
�  *�  *�  *�� +�� �  
�  *(  *
  (
  ��    ����������������  ��  ?�  �  �� ?�� ��  ��  ?� �?� ���?      �   �   �  
�  *�  ��  ��  ��  �  
�  *(  �( �   �(     ����������������  ��  ?�  ?�  ?�  ��  ��  ��  ���� ��?��      �   �   �  
�  *�  *�  *�  �  �   �  �  �  �   �     �������������� ��  ?�  ?�  ?�� ������ ��� ?�� ������ ����      �   �   �  
�  �� ������
��,
�  
*  

� (� ( � (      �������������  ��  ?�  �  �   �  ��� ?�� � �� �� �����     �  �   �  ?�  �� ������ ��  �  �  ?<  <<  �?  �?     �������������  ��  ?�  �  �  ?�  ��� ��  ��  ��  ?�  ?���     �  �   �  ?�  �� ������ ��� �  �  ?<  <<  �  �      �������������  ��  ?�  �  �  �  ?�� ��  ��  ��  ?� �����     �  �   �  ?�  �� ������ ��  �  �  ?<  <<  �?  �?     �������������  ��  ?�  �  �  ?�  ��� ��  ��  ��  ?�  ?���     �  �   �  ?�  �� ��������  �  ?�  <�  <<  �?   ?     �������������  ��  ?�  �  �  ?�  �� ��  ��  ��  ?� ?����     �  �   �  *�  �� ����� ��  
�  
�  *(  ((  �*  �*     �������������  ��  ?�  �  �  ?�  ��� ��  ��  ��  ?�  ?���     �  �   �  *�  �� ����� ��� 
�  
�  *(  ((  �
  �      �������������  ��  ?�  �  �  �  ?�� ��  ��  ��  ?� �����     �  �   �  *�  �� ����� ��  
�  
�  *(  ((  �*  �*     �������������  ��  ?�  �  �  ?�  ��� ��  ��  ��  ?�  ?���     �  �   �  *�  �� �������  
�  *�  (�  ((  �*   *     �������������  ��  ?�  �  �  ?�  �� ��  ��  ��  ?� ?����                                                                                                                                    Z\^`bdfhjlnprtvxz|~���������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLZ\^`bdfhjlnprtvxz|~���������������������������������������������������� 					
		


 
"
$
&
(
*
,
.
0
2
4
6
8
:
<
>
@
B
D
F
H
J
L
Z\^`bdfhjlnprtvxz|~���������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLZ\^`bdfhjlnprtvxz|~���������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLZ\^`bdfhjlnprtvxz|~�������         
                                                                                                    tuvwx                                                                                                          ���                          