��N�  r   
                      P �                         h � � (
 h � � (�j � � *
 j ����*@l � � ,
 lP� , n � � .
Pn0���@p � ��0
�p�����0�r � ��2
�r0����2`t � � t@����4�v � � 6
�v�����6px � � 8
 x��p�`8�z � � :
 z�����:p| � � <
 |���<`~ � � >
 ����>p� �  	 @
 � �� @@� � 	 B
 � � �B`� � 	 D
 � � D@� . 4
�0~�                 � � � �𠠠���  ����� ������ �  � ����� ���� � 2,���#���#�����#�;/�(����������      �� ����   � ��� �� ��� �	8 � � �� � ����    ��   ���  ��� �   
   ���� 
���    
��� ���� �� ���ʯ���
/��Ԡ�ST�P �?����@ ��� � �  � � � � 2����     
 
 
 
�  
��
� ���>P��
� �
 ����   �U�  �!P      
     ��  ���  
 
 
 ����        �� � �
 
� �     �   �����,�:�����0L���       ?     < � ��   ���      �
�    ��
� �#�
?O<
�/���0
�wpW      0 ?     � �  
    ���       
    ���
�,�#�
;?O<
�-���0
�wpW        ?   0; �  3
    ���       
     ��
�(�#�
��O<
�-���0
�2wpW 