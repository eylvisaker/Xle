�6287	 ��;|�      � D                      �      �   � �     � @     @ �   @                                @                             �               �                  
�     @   �  �     ��      �     @ � 
����     @        *ઠ�             ��

�             
�� ���           P�     �         Z ���        A   ^  ��  �       � +
�           UU`             UU�  
���@          �U�  ���         U�  @ ���           UT   �� � �      P��  �
�         ��P?�  ��     �   ��U��
���    �     ?�� >�����    @    �����������        ��������      �����껻���        �������       ꪪ������� ��     �� /���
����  @    �� ���������  �   �� ������  @   �  �
��������     ��  .���������      �� ���?�������      ��
�����������         �����������      
�
�  �����  �   �����   �����     �����    ���� @     
1�J8    ?���      ʆ�*     ��    �Ҫ��0    ��      p **��   ��         �     ��     @     �   ��        @�p     ��      B    `   �   �              �               �     @                   @       @                             �      �          �       �     � � � �     � @                     �                                      @                                                                          �   �  � ` )                                    @   �             ��@     �*��   �     �"� �     ��
      
��%     
� E    @  +�U       *�  u  �  ��� U     @� ��     ��/�S�    ������   *������     ��ȯ���    ��;��*�  ������   ����. B�  ?����
�   >�����   ��� *��    ��  **   �� @ !$�    ?�  �*���  >�  B� 4  ��       �@       �  @�                                @   @                 @ � @     � � �         �  �        @                   *  @  ��   �     E��  @ T :   t .�  �"�@ ?��:�   �����   �����@����   (*���� 8����  �  �� ��i��� (0 � �@ �       �    @  @               �     0     �B  �    � 
�  �+�   .P�� � P �H  �>o @ �������� ��� @��"� � 	�� ,�  0 B     �  @  �     �         @    
� `�@�@(�� ��+�������    @ �� @	 ��;|�      � D                                                           � � @   @ � @                 � �                         @      @                                                                       @ @ @                           �       �     �            @ @   @            �                     @          �                 @                     @ @   @        0       @    �   �     �      @ @   @�               �             �    @           � �     �        � � �           ��  �  @ @     � 2   >          
� �`  �       @ @��s� �  �       � ����&c��     �  � .�O�	�       � 
�Ϻ{�          
� w>�ߨ �       
� ��� fw`�  �  �  ��wwt��� �     � ������&wv ��   �    *gwwO������    @�  
�����wvo��   � gwwO���ڠ <   �  ����fwwv @�   /�  7wwwp���  � @ /� ������&www  �   *��%wwwwO������  
�������Ϯ&wwwp �  ��gwvwwN
���� ?�    *��������fgvwwo�� � 
�wwgwwO����ݙ��     ��ݝ��Ϯ&vwgwvj�    gwgvwvN�)ݝ��٘    ������  fgvwgv�    &gvvvv`��m���ߘ    ����ٙ����vvwvf    f�fvwd��f�%��ٙ�� 	����٘����vvfffd   f fvc�@o��ٙ 	�   �	 	�������fe  e@  @fef?o��A��	��   ���P����"/�f`o��`   ������H��@����   ��ff��"/�d ���  ��� �Ȉ�`	�  �    � �"/� f  @�  @ ����@H� �  oə   g��f�  ߐ     	���d ���	�     ���� f	�`�    	��f ` ) �      �     �   �                      @�      ��    �  @     �   @      �           �   �     @    @    �          �               @ �     �  �        �      ��      @�  �   � �� < �    �� �   �  *s�_�� @   	�ៀ0  �7B
v <     ���ᝃ�    �ws�w� � � -��)�� � � wws�wx  ���Ӊ�� ���ww|&ww  +���Ӊ����  
gvw{�g{w� ����!�ݝh vfwO�ggw@  ���o��� fff佋�fff � ��gf�	� 	�a���`&`  ��A�r'��� f� d+�� �   ~	��'�@�ـ  @ ��`FB@��      @   �                         @     �   @              �    ���  @�0   �   ��8  ���� ��܉��  ��w'_� �܉� �ww&w ���܉��� �ww&w_����܉٘ fgt'vf@  ��љ���&<�d& , ���	 ^A���    @�0  �      �                       � � #�   ã  � �@0&��  .tɎ 	܆z ,7w)�0�܆v�vw)��	��f`$cƘA�1B@�M��� x          @�    �    3��;� ���0v��.lfx	��F�$	 @  �	 ��;|�      � D       �                                  P  @��  �        U     ?T        @ TP    UUP  @     @P T   P �         P   T  ?@        T   @  �@ �    P     �@       P  �@ �       @   T  �    �      P S�   �       U@�     �    @   T�  �  �    �  U�    @ �  @  �w �@�T    ? P X�� @�U@    ��T  �#p C�P    �� U  4�� �@       ?  �g@U� �� �   @ ?� T��� �����P � @?�< ?  < ���P | C� <      ?��T�  U?�@< �    �?�UE� T��@�  � ��UW�AU_�P �� @0?�? �S�UU�� T  �   ����O�T���   ?    � �?U_�U�T P �  P �?W��UUUU@ U�  UU 1U�U��UUUUT �  !TU@UUW�U?�UUTU�� �@UUU�U��UUC��   US�U_��UU�_�U    ��U5������T  @   �UW��U���U @  P  �UUwUUO� <@@    ��]UUT  P@�  ��UU��UU   UU     ?��U_��U@ � P   P��UO�?�P      @   �UU?��T          �UP��� U  @   �?UU� ��P �      _U@?�  � U@  �   UUT �   �UUT      UUUP�  ��  UUP    UUU� @�   UU@ � T@ �� � UP  P�  ?� �     T   U@? �?   � �  U U   ?   ?�   U  P� ?   �      @ �?    �   �  �@@? �  ?�     @ < �   � �   @   �     �<�  @P   �   @ ?�   P <   <  UP   �T  T <    QT  @ P   U < @U T  �U@  P   �     T     T<   �   @  S     � ��<  P  U         ��  U UT�?  P �   ��  UU@ ���U     �   U   ? �T      � �     ` )    �� P    T?       @  P @ @�  �    �       @   �     �   T        �  <P    �   0PP �   �P2 P� � �@x� @  �@@@    �B� <   � 0P ��   �<U�<�0 U�P���@0�S��C�    < P���??   AT��S��P  �UU}UU U  ��\QUUP @ PS���T�T@!A@?�U<  U W�O��@  T C��P� @   ��U5P� @T? <UU   U@? T@ @ ��T �P @� @ @� <  �<P @ � �< �P@?�  @ S�    @� �PP T @@ �<  <U � P0� P �  T  �  �P @   �  @P@    @C  �   @�  � T�� 0 �@<R �P:A=   0| <  <��}T� �}_�ÀP3Q}}E<UuUA@U7]s�R�H�=_  <S�T!@]C�  �T P�<A 0�� 00�?  �<@�R @�@@��A@� 0P0   @�@ �P    0P� �1@0� ��i0  �� 21_� �_ ?W]W�@|U�TM_ @s�� T��U �@<01P�<�� 00 P�0@<A �0# �Q    B  ��� �dЃ�� =�sSW�=��W=B�<����@	 ��;|�      � D                              �   �      �@ �   � @ � @                        DD                             D@                          A      D       �    �     �          � @   @ � �   �                       @                             @    @   �        �     �          @    D      @               �       D@     D@   @                   �          D                       @        @          ��        @@  
 (    D @       �            @ � �             �  �             ?�  �   @          � �          @  ��+�    @ �         ���          A     ��     D  @                      D           @                         @          D@                      @         @@                 �     � @        D    @                     @                                  D@         DD@                    @@           D                                                                       @                     ��D             @                       D                                �                  �                      @                @D@@                      @      @ D@     �    @@ �    D@         �    �   @  @  D �        D  �        @   �  @DD      @              @` )                       @  �    Q   @       @�       D    B     @ ��     @        @    @                 @            D �  D              @    @(2     � �     � �      ��      �             @                @   D             @   �              D         @          @                   D        D                  @            @    �       @DD D  D       D@  �D      �   @   @ @         @ � �       @      � @ �    @      (  @  B�� � � @ ��    <  B             @             �      @           �@    �    D@DB    �� � � 0  �        @ @   @   @� D   @ ���  @��  . �@    @    @ @   �    B    @    DB DDP �    �   �@ ! @�  @ @�0�H  �  B  �D @   �	 ��;|�      � D   @                    �  @         �      @       �  @                         @                
 
�             � *���              ����              ���      �@      /���       �        ?����    �        ������             ������           � ����            U���@    @�      UU���P            
 D���P    @     � 
   ���    �     @ � 
UDO�     @     @  ���@       �      GD��P          ���             � DO�T@  �            _�Q�       @@ @   ��D��             ���@         �TDJ��P          �����    @        
�_���@           ��      � �   � D��D��             
��P           ��DD��P     �   �  
�����      @  @ �����O            � �Z���    �     @
�DD�D��            ���P            �DJ��             
�����P �  A  @    *����@             ��ڤD@          ����         @  �DDD��              ����        ������      � D�  
������       �� �����D    @   ����M�����   �  _�_���<u���TO�     @��5�DD��Q�      �G����DEUDD�@ @   ���_�O�*�     D������DD��@�    ��QO������      OQ_���������     �T_O���ڡ�   � OG�QQ�DU�TDJ@�    @����!Q��      �DGuE���DDDJ��      U��J����     D]E��M���TJ@     Q_�աwQ��@      D_����DD��� @       E_������D�    �  @ �����U�       
��J�O�DDD
�     �  �   � �  �` )               �               @  �        ��  �    @ ��     � �4��       �?��     ��A�     ��T�    ��� �      �G    �  O�    ��   �D      ���       ��       �F� � �  ��
      ѯD(      ��  @@  ���      ���@(  @  ��� �  �    �F       ���    � �iG      � @     ���� @    ���@� � ��A���    =�4D}G@   �DH�?���� �Q�}?���  6���=�P   EUT�q]�  *(��OL@  !�D���  � *DS�TD   +�D���A     !?��
�   
 D@� * @� @  � @        ���   ���     ��   D�� � �B/�     ��  @  �   �0   
Ҽ � (�    ��  �����   
F�   	�� �   (XD  k   7@
��@  qs��B �Mr�[  |v)@�Q=UFB �SN�V�@ G�=�   ���F� ��(0           � � �   �X x   = � !O�@  � @ =�    [ր  o  �h  i  @��@ ����E-4� U\EL 
D��
��  H
       � @�  �@�  p  ��    �� %@ ?��G'�]d�s%((U 	 ��;|�      � D       �    �           �   �   p         �   �  4 @        � ��   =         @ �  �   }         �� �  ?�           ���
����         �������@   �     ���*��              �� ��@           @  ����
    @      ��
��� (          (
� * *�         @  *��P�
��    �     (��   ���         ���ꊪ��    A        "� ( �(          @ @"��(
�             �����              �����   �     @  �(��(�        @   
��
� �"�           �����"
����         
�*� � *�"��   �   *ꪪ�*������      ���"��"*���       ������ �����    �����""""���      �
���ꪈ��������     
������""������  �  *����+������*��      *�*������������    *�*�������*����  @   ��*��*��������     ��*������������     ���������������      ���������������     �������ꪢ��*�*      ���������ꪨ���     ���������������      ��������������� @  *��*��ꪪ�ꊪ��      *��*����ꪪ����      +����������*�*�      *��������ꈪ���   @*��*�*��������     
��������������     
���"*����"�*��     
������������� �@   ���"(��"���      *��������*�      �*� """ "��(        ��� ������     ���"    " ����       *����  �����      @*��"  " ���  �    
���     *� @      ��   " *�       ����   �+�        ��"   " *�       ����   �*�      @  �"   " .��  �    
���    �*��    �         �  �     *
��       �*
�    
*���     ��*�     
*
��      ��*�    <4�    <�� ` )   �  ��        0     <   4    �@�      ����@  �    �
�       
*�     
���      �� �     �����    @ �#��� � @    �*�      �� ��     ���* @ ��*���   
���"�    "��� ���    *��"���   �*�ꪪ�� @  �**�.����  �*ꊊ���� �*��:���� ���������  ꋢ�*ꢪ�  ����*���� �������
��   ��.�*�*��  ��*�*���   *������ � .�*� ��    
� �����    *   �   �� �*�   
�"  +�    �    *�@  �" "*�     ��  *� � �"  " �    *
   ��   ��    0� 0�        @      0  0   <@<    �+�   ���   �� � ���    (
   
""(  �.� :����  
���� 
*����  *(���� �"*�(��  :�**�� *����� .��(��  *��**� �
�(�*� (
 *   �� �� � 

�  �� �  �
���� 30  �   ��0  �    @ � �   �/  B "�  $   
( �  ��  
��� (�* "���  �*��� �*������*  �:"+ *�� " �  * � 
 � �
 �  "  �0� @      ��0 
� ��  �  �
�����** ���B��� � � �� � �3 ��