�Y�  �HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHg���HHHHg���HGGGGGGGGGGGGGGHHHh���HGGGGGGGGGGGGGG HH::::::::::Hh���HGGGGGGGGGGGGGG()HH:::::::::: ���������Hh���HGGGGGGGGGGGGGG!)HH::::::::::.0�g�������Hh���H<<<<<<<<<<<<<<!)HH::::::::::/1�h�������Hg���H<<<<<<<<<<<<<<!)HH:::::::::: �g�������Hh���H<<<<<<<<<<<<<<()HH;;;;;;;;;; �h�������Hh���H<<<<<<<<<<<<<< HH;;;;;;;;;; �h�������Hh���H              HH;;;;;;;;;; �h�������Hg���HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH;;;;;;;;;; �h�������Hg������������������������HHg�������HHH;;;;;;;;;; �g�������Hg������������������������HHg�������HHH  (   (   �g�������Hg������������������������HHg�������HHH***�h�������HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH�h�������HH�h�������HH�g�������HH�h�������������ATTTTTTTTTT@HH�h�������������SATTTTTTTT@S ***HHHHHHHHHHHHHHHH�g�������������)SSATTTTTT@SS )""")HHh������������H�h�������������)#SSSATTTT@SSS.075555555555555554HHh������������H�h�������������)#SSSSATT@SSSS/1-755555555555554- HHh��HHHHHHHHHHH��������h������)#SSSSDBBESSSS --7555555555554-- HHh��HHH���h������)SSSDBBBBESSS ---75555555554--- HHg��H�h������SSDBBBBBBESS ----755555554---- HHg��H�h������SDBBBBBBBBES ----822222229---- HHh��H�g������DBBBBBBBBBBE ---82222222229--- HHg��H��������������g������            --8222222222229-- HHh��H�������������(�HHHHHH�-822222222222229- HHg��H�������������%+82222222222222229 HHh��H�������������%+     (   (       HHg��H�������������%+***HHh��H�������������(HHHHHHHHHHHHHHHHHHHh��H������������� Hg��������������HHHh��H������������� Hg��������������HHHh��H  (%%%(      Hh��������������HHHh��HHg��������������HHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH;%   99;IKM?75++AKMEB=�����%	&&%$"%%$�����
 9� '� GtC t%" "
�����������  o� ����  o� � �f�  -� ��f���o� ������o� � ���  -� ����  o� �� ��  o     �����   ����+���������������o � - ���-  ��o��- ���-� ��o��- �---�  �o �--ȗ����  �o����       �o           ����������������(GGGGGGGGGGGGG ��   o�  GG   � �o�� G  � � �oo� f  � � ��o��f    �  �o��GG�� �� �o� GG��� � ��� GG��        GGGGGGGGGGGGG�;[[[[[[[[[[[   [[[[o �-�          [[o�-�     ����[[o�-�     �-���[[o��-�     �-���[[ ��-�   ���-��[[ ��-�   �---� �[[ ����   ������[[               [[[[[[[[   [[[[[[[�	______________�β�      __�ε������  _��ddddd��  _���������  _ ��������� __           _____   ______�������    �  ����   ��� ͧ          ͧ������    ͧ������     �   ��� �   ���������������������4��4�  �4��4�  �4444�   �����                  ����������D
�����������OOO     ��O ��� ��O���4� ��Oȳ�4� ��O ȵ�4� ��444444� � ������� �         � ������� ��444444� ��������� ����    �� OOOOO  ������������-----� ---------�  \\  �-ȳ���  -ooooooo-�  \\  �-ȵ���� -o�

�

-�   \  �-���o- ��ɳ��-�      �-ooooooo-�  ɵ��-�      �--------- �------�  \   ���������  ��������  \\                       \\\\\\\\\\\\\\\\\\\\\\\\\\�[[[[[[[[[[  [[�����������[[��������� �[[ � � � �� � [        ��� [� � � � ��� [         ��[[[[[[[[[[[[[[�A              ( ( � � � r  L A S T   C H A N C E  P I R A T E ' S   T R E A S U R E  C A P T A I N ' S   S H O P  D E A D L Y ' S  T R E A S U R E   C O V E  T H E   S U R G E R Y         