�Y�  �UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU}UUc����������dU*+�c��������da 33334444*$��c������daa 00000000000000000}33334444 nimnm*$��daaaaaabaa 00000000000000000 U33334444 ijjijm�daaaaaaaaba *+00000000000000000 UU33334444(*pil pil�daaaaaaaaaab *$00000000000000000 U33334444 *              *$///////////////// U33334444 **$///////////////// U33334444 **+///////////////// U33334444(*///////////////// U33334444 LPPPPPPPPM     (   (       U        PLPPPPPPM�****+UUPPLPPPPM�� UPPPLPPM��� 			jkiiijkjjkijijjkkkiikkU����������������	PPPPPPLM���� 			krqutqrsttrrui		iikjjjkiU�>>>>>>>>>>>>>>�+PPPPMN���� 			irtruqqrtrrtqi		UU�>>>>>�����>>>>�+#PPPM��N��� 			ktqsstsqssuqti		U�>>>>>�����>>>>�+#PPM����N�� 			ijiijijkkikiii		U�>>>>>�����>>>>�KKPM������N� 				












		UU�>>>>>>>>>>>>>>�M���LPLPLP 							**@@@@@@@@@@@U����������������PLPLPL 							*!@@@@@@@@@@@ U		














PLPLPLP PPPPPM	*!@@@@@@@@@@@ U	kkik	P       LPPPM� ����*!@@@@@@@@@@@ UU	kjjjPPLPM��PPLPM�� ����**@@@@@@@@@@@ U	kj
]]]]]]]]]]PPPM���PPPM��� ����AAAAAAAAAAA UU	kk	]]]]]]]]]](*nimPPM�N��PPM�N�� AAAAAAAAAAA(*U	ki	]]]]]]]]]] *oijjPM���N�PM���N� ****AAAAAAAAAAA *UU	ki	]]]]]]]]]] *pil M�����NM�����N *""*AAAAAAAAAAA *U	jk	]]]]]]]]]] *               WWWWXXXXAAAAAAAAAAA(*U	jk	**^^^^^^^^^^(*WWWWXXXX            U	

	*!^^^^^^^^^^ **WWWWXXXX *!^^^^^^^^^^ *!WWWWXXXX UU*!^^^^^^^^^^ *!WWWWXXXX nimnimU				iikikki^^^^^^^^^^ *!WWWWXXXX ojiijijU				






          iiiikkikkijk+WWWWXXXX pjl pjl UU												kiikkijkikjjWWWWXXXX   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUK>BGLLL2L!H�������������$#	�������������	, $x 6� ?� P!((3"�7�?�K������������    �������Ա������Ա�       �����   ���O4�  ���4O� ����������%�������������  � �����ר   � �����ר   �   ���ר   �   ���ר�������������7������������������    ��4�       ��  �ȵ�4�       �   �4444� ����� �   ������ �444� �          �4�����         �4�����������   �������� 
����������� ������ �����   ��̵����� ��444444� � ������� �         �         ��        ������    ��$�    ��#��    ���������       �4��ɱ������� �4�� ��4O4O4� �4� O��  ��O� ���O��  ��4      O����������������
�����������OO�    ��O����   �O��4�   �O��4�   �44444�  � ������  �         �         ������������4���  ����    � ��    Θ�   ����   β���   ε� ��  �11>��  Ξ����@�����������        ���        ���  ���   ���� �4�   ���� �4�     ����4�     ����4�      �  4�      ������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                A       
         � x x d  U R B A N   C R U N C H  S T R E E T   S H O P 
 C I T Y   S T E E L      T H E   G E N T L E   T O U C H  H O N E S T   A B E ' S  S H A D Y   S A R A H ' S    D E N   O '   D E L I G H T 