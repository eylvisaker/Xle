��N 7  � A   
                                                � � ���p(�j *
 j ����� ,
 l`.
 p � 0
 p � � ��2
�� �@��4
 t0� v �6
�� 6 � 8
 x � � 8 z � � | � <
 � � � >
 ~ � > �  	 @
 � �P  @ � B
 � � B � h`(
�hP����*�l@�p�p��,�np� ��n@��� .����0�r`r��p2ptp��4��pv��`x��@��:
�z0�P:��@|�<@~����p� �0	`���	�D
��p��0D�                &`                            ?�  ?���;������
�  5���T��u]UP���������u������    � ��  � �������W��w��������  ������� ��������U�UU_�]UWUUUfdf`f@d ����� �  �?��� ��?�����?�� ���?�� 	���������������������fff��������� � fpfd� ������                                              0                       0      0                 0                0                   0      �U]�UUU��uUUUU��U@UJ_���U@U�����@ _���u _�W�U �@���     �       ������ �����     ���� �  ��
� �    ����  � ���                                               0                       0      0                 0                0                0  0      �U]�UUU��uUUUU��U@UO_���U@U�����@ ^���u ^�V�U �@���     �       ����� �����     ��� �  ��� �    ����  � ��                                               0                       0      0                 0                 0                0  0      �U]�UUUo�uUUUU��U@UO^���U@U�����@ _�ֿu _�V�U �@���     �       ������ �����     ���� �  ��� �    ����  � ����