���$ G  G	 Q  Q c  c	 {  { �  � �  � �  �  $ �       '  ' 3  3
 A  A
 U  U i  i  � o �  � �  � �  � �  � �  � �  � �  �   �       #  # )  ) /  / 5  5 ;  ;  [ ? [  [ ]  ] _  _ a  a c  c e  e g  g  y i@�t �$B)                                                                                                                                                                                                                                                                                                                                                                                                         �$                    � �  � �   �     #   - #  5 -  = 5  C =  G Cf	�	�	&
	f	�	�	&	f	�	�	���"		�F
"	����"	F��"	����	,
	l	�	�	,	l	 	�@
����"	 �@���0
	p	�	�	0	<
�|"	���"	<�r2	�2	�	22	zB	�"	�B	:�t2	�2	�2	xB	�B	6"v�xzt�t�~�n�r�z�x�p�v�|�t�:p�x�|�~�v�n���r�4z�~R	xr	z�	r�	pr	n�	tr	vb	|r	|�
pb
x�
v�
rr
z�
t�
��r0B��2R��z26r8btx��v"��:�p�4b��46t�x�v�8�r�2"�R,
bl����b,�lb�b���B���2���"���"������"������������� 	�@
r���� r@��r�r r�R�2�B�r�b�b�R�b�2�R�B�2�"�B��	��	��	��	��	��	��	��
��
��
��
6�
4�
8�
��
2�
:�������r�b�B����R���B�R�2�20
bp�����0�p����"2
����4
����6
����8
����B:
����R<
r|�����<�|����b���r��2�"����b�r�����
�
��	�xBvB�"tB�2�"��xv�t��t�v��rx����b2
2r���r2rr�4
t�t�6
�v�v�8
�x�x�:
Bz"�R�b:Rzbx�v�v�t�x�x�v�t�xB
v2
t"
�R�r�bv�t�x�t�v�r�����2�4
�t�6
�v�8
�x�z��:6�6B6�6R
6
�626��"�24B�R6��b�r8�fjf��fnn���隚���ff���f��������jf��f�f��������jff��nf����������f��f�f���������jjf�fff��������       
    �� 
    ��  ����  
         ��           
  ��(       �     ���    
       
      ��(             ��             ��� �   � �      �       �       �     ��       � �  � ��         
    ��         �         ��   ��     � �      �              �        *�  f�jjf�f���������    � j�    � ��      ��      ��
��f����)�������     ��     
f�"&&&fff ��������"""&jf  ������  &"�&�� ����������j�fjf���������    ��ff    ����
f*f�ff�	�������` j f��"� ����HH 
 �f��" )����HH    f��"  ����HHff��"""���������jfjff�j�����"���j�fjfjh	���"!����  jjjf  ��""��  ��������"""""  � ��    
           *     
 �  **� � 
�� �     ��    ��        �� * �� � 
      � �     � �   � �     �     �� 
��   ���    ��  ��    ��    
�� ��  ( ��        
     
     �   ��   
�   �
���  �* ��  ��  ��      ��  � ���  
� ���     
 �     (      ����             EU  Q@TP P  UETAPPEUUQTUUU PPQEPPEAEQQTQTUUU PDUPDPEUP    UUU  PQP      P       P   �         E  TP  PQQP  UE    UT@@@TQ   @  U Q  @      P      PPEU   EP    A@P    A             A                   Q   ���     @    P    �   @       �z p�

��Р 
� �  *�    �
�    � 
��   ����   
  �               �            �
Z�P*
 ��R� 
�     �  �  
 * �    *��   � �� (   P�
 �  �R
�       
              �    
�         H�   @��            ��  �      @ � �� 
J            ������w�������U��������������UU      ��    �@UU      ��    ��UU      _�    ���U             �U U��������UU����UU� � � � U � � U  � W     �     ����    ��UU    � �     � P            _  �   �      ��     UU      ��    UP_�         UU��  ����                  P  � � � 
 ��� �  ��������������%�����������������������𪪪������������������� Z � � � � � � ���UU��������������UU��������������UU�
����
�
�UU������������      �P    U ��      ��    UU��      Z�    UU��             Z*j*j j  *j
j        �%U  	Uj*j    ��UU  UU���
    �@UP  U �P��������  ����    �
����  �
��        UU�� j��*   * * *  * * 
  ����������������
�𪪪������������������������ � � � � � � �      )     *  UU��UU  j�����  UT��UU  ������    � T   @ � �   
 
    
   ��j�j�  UUj�j�  � � �   U � �     UU��UU  �����
��<  ��� ��0 ���< �< <   <��0��<��0 <0�?�������<�0� ����� � ��������� � � � 0 � � �  � � 3 � 3 � 3 ��0� � ?��?����<30<<?�3� �?�  ��<0� � � � � � 3 � �  �  � 3 3 3 < �                      ��    ����  ������  �������?<<�<�3��� �<<3�����00������<���<<<�<3����3�������<���<?<�<<��� �����3���0���???���<� 3�0���00?<�����0?0�����3� <��0 � < � �  � < �   � 3 �  0 ����<� �<     � < � � 0 � 0 �  � � � 3  3 <�<�<�<0� �3�0� <<�  0������??�3��0�����<<�<<<� � �������3�<<<? < 3??�?����������0�������????3?3? �  �   3 3 3  �  �  3 3 3�  � � 0 � 0 � �  � � 3 3  0     ����  ���������  � �  ��<�<������<<00���3?�3���?3�<���0��<���3���������<�����������������������<��?���<���?���?���?���?���?���?����<�0��<<��<<���< � < � 0 � < � < � ����0 � �������0  <<���  <?�?<<��<<0�� < � <   � < � < ����  3����    ����    ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              