��N�   x   
                       P �                         h��@�@(
`h@�@��(�j@�p��*
@j@�p�@*�l��@�@,
@l@�@�@,�n��@�p.
@n����`.�p��@�@0
�p�����0�r��P��2
Pr0�0��2Pt@�@��4
@t@�@��4�v�� �P6
0v0�`��6Px��`� 8
�x�� ��8Pz��@�:
�z�����:�|@�P�@<
p|p����<�~��@�@>
�~@���`>��`�p 	@@
@�P�@ @@����@	`B
@�p�@�B��@�@	pD
@�@�@@D�                PPPPPPPPTDTD    ffffffff�������   D   @@D D    U@D@PP@@Q  PP    D �   ffD   	���   fd&f  	����� fff&fF	�������             	�
P
P ZPZ�  ��  
P
PPZPZ�  ��� @@@@DD       D      @ @             DD  DD      DD  PPP     P PP  DD@     D @                    @@ TPD   Q  &ffffbbf��������ffbffbFf�������    �� �    ��      �  P    U�      � P    U�     ��     UP     �P    �U      �P   �P      �P    �P   DDDD    D@ DD    DDD@    EDTDQ    U__
Z�  U  T@DDQ    D@ D  