�y+N
   x   
 0                      � ����                  h@�P�`(
0h�� � ( jp����*
Pj�� � * l�����,
 l�� � , n�����.
pn�� � . p � � 0
�p�� � 0 r0�0�2
@r0��� 2 t0�0�04
0t0��� 4 v0�0�06
0v0�0� 6x0�0�08
0x �0�@8 z0�0��:
Pzp����:�|`���<
`|�����<�~0�0��>
�~� �0>@�0�0 	0@
 �P�` p@��0�0	0B
0�0�� B��0�0	0D
0�0���D                 DDDDDDDDDDDDDDDDDDDDDDD@ D D DDDD DDD    �    
@            P @ U  P  DDD D�D   D   @@P�  @ �
�   Z��  P @          P  �   ?��  �<�DD DD D    DDDD D     DzDzDzDz::::      �       ��D D         DD  @               DDD~DzDz:::: 8   � �    � � �  # � 0� DDDD           @P  @                @      D     P     DDP   DD D          DDDDD   DDDDDD   D   @    DDN � ��8 � ����������������D�����OU@UOUOZUUU�DUTDTD�"QQY��L*���� �U""�L*Oʨ�0�O
O��UUS _
�_U
��?��ߪ���������U?�����?����?���������������O����5T�����PU������  _��_�  DDDDDDD��DDD@@      @"" ""*"���������"*�
*R�����B�Ԩ�
P����������������� �����U DDDDD D����" """"""��������""�"
"P"��(�B��   P    @ T U@DDD$D" ����"""     ��      DDDD@    ��* " � * ������� �TE�D�uUU]UՉUDDDDDDTD QDzDzD@G]: ��DDDDTDDDQQ               """""""*��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              