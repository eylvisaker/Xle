��NZ   x   
                       P �                         h � � (
 h��p� ( j � �*
0j@�P� * l ��� ,
 l�� � , n ��� .
@nP�`� .�p ��� 0
 p���� 0 r ��� 2
 r � ��20t��p��4
�t����04�v��`�@6
@v@�P��6�x�����8
�x����8�z ��� :
 z � ��:| ��� <
 |��p� <0~ ���>
0~@�P� >�� �� 	 @
 ���   @ � � 	 B
@� �` B � � 	 D
 ���� D                 ��  �������j�j  ��������`���� ��� ������O?����_�?�� ��� �����ꪪ �� 
�*��� ���  �ꪪ��:�����             :      �     � �           ��      � �  �����UUUUU@UUUUU@UUUUUUPUUPPUUPUUU

U
�U�U ��  ����n���  ��  ������  ��  �����着��  ����	�	;	 9U
U
U
U�UUU�U ����    ��      ��*�    ��      ����    ��             �                 �  પ  ����������      ����  ���  ��  ����������  ����������������
�
�
�
�
�
�
�
�����
����  �    � �  �� � � �  � 
 
    � � � � � � � �  
 
 
 
    ����    ��