��N    x   
                         @                         h�����(
�h���� ( j�����*
�j�� � * l�����,
l � � , n����@.
 n�� � . p����P0
0p`��� 0 r����`2
prp��� 2 t�����4
�t���� 4 v�����6
�v���� 6�x�����8
�x�� � 8 z�����:
�z � �P: |�����<
 | � � <�~�����>
�~@�`�0> ��� 	 @
 �P�p @@ ����	 B
 �����B �0� 	 D
 � �  D                                             @     A   ���������������������������������������������������������*����������������������������0�������  ��������"""""""";�� �  ��   ���     "       �������
������  � ��  � �   
���
 �� ��
��� ���
 �
�� �

� ���������
 *
���� ���* �*������
������� 
�����������������������������������������������������"**""*  ���     � �     ��������������પ���   ��� �   ��� � � � � �   ������� """""   ����    ""      ���             ������� """"" "                 ��������""""" "     � E   4UU  U�QU� UWUQUU Q T Q PUUUUUEU@P   EUTUUUU    @                    � � � �                          � �         �������("*�"������������""*""**"��������"""""**"