�Y�  �HHHHHHHHHHHHHHHHHK������������HIIIIIIIIIIIIIIIIIIIIIIIIIIIHh���������HHHHHHHHHHHH������������ Kg�����������H++jkjkjkjkjkjkjkjkjkjkj Kg���������HvvvvvvHH������������(++%jkjkjkjkjkjkjkjkjkjkj ++vvvvvvHH������������!++%jkjkjkjkjkjkjkjkjkjkj +%vvvvvvHH������������!++%jkjkjkjkjkjkjkjkjkjkj +%vvvvvvHH������������!+++jkjkjkjkjkjkjkjkjkjkj +%vvvvvvHH������������(+KhmnmmmnnnnmmH      (    (         KhmnmnmmnmnH++vvvvvvHH������������ Kh�����������H++++++Kg���������HvvvvvvHH������������ Kh�����������HKg���������HvvvvvvHH������������ Kg���������������������������������Hg���������H++vvvvvvHH     (   (   Kh������������mmmmnmnnnnhmnmnnmmmnmnn���������H+%vvvvvvHH+++++Kg����������������������h���������������������H+%vvvvvxHHKg����������������������g���������������������H+%vvvvxwHHHHHHHHHHHHHg����������������������g���������������������H++vvvxwwH�mnmhnnnmmmnm����������������������h�������������HvvxwwwH����g������������������������������g�������lllllvxwwwwH����g�������������������JIIIIIIIIIIJ�������liiil�xwwwwwH����g�������������������HKg������liiil�(   (H����g�������������������HKg������lllll�+++++H����g�������������������H:::::::::Kg������     g�����HH��JHHHHHHHHHJ�����������H++::::::::: Kh������g�����HHHHH��HKh����������H+%::::::::: Kg�������mnnmnmnn������mhmm��H+++++Kh����������H+%::::::::: Kg����������������������g����H+%%%+Kh����������H+%;;;;;;;;; Kh����������������������g����rllllllllllqKg����������H++;;;;;;;;; Kg����������������������g����prllllllllqp Kg����������H;;;;;;;;; Kh����������������������g����pprllllllqpp Kh����������H::::::::: Kh�������������MGGGGGGNHHJ���ppprllllqppp Kh����������H++:::::::::(+Kg���������HHHH<MGGGGN< +++++Hg��pppprllqpppp(++%::::::::: +++<<MGGN<< +%%%+Hg��ppppprqppppp!++%;;;;;;;;; ++%<<<MN<<u<<<<<<uHg��pppppstppppp!++%;;;;;;;;; ++%<<<><<u<<<<<<u< Hg��ppppsootpppp!+++;;;;;;;;;(++%<<<><u<<<<<<u<< Hh��pppsooootppp(+         ++<<<>u<<<<<<u<<< Hh��ppsooooootpp Hgnnmnnmnmmnm�����������������nmmnmnnmmmH<<<POOOOOOOQ<<< Hg��psooooooootp Hh�����������mmmmnnmnnmmmmnnmmn���������H<<POOOOOOOOOQ<< Hh��soooooooooot HHHHg��������������������������������������H<POOOOOOOOOOOQ< Hh��mnnnmnnmnnnnmnnmnm��������������������������������������HPOOOOOOOOOOOOOQ Hg����������������������������������������������������������H               Hh����������������������������������������������������������HHHHHHHHHHHHHHHHHHHHHg�����������������������������������������������������������mnmnmnmmnmmnmnmmmmmn @=?BM;<, 
8G���������������$"!���������������
8 8 !� +� HHL��!!+=�I�[[[[[[[[[[[[[o        [[o����     [o� -�     [o� -�     [o��-�    [[o��-�    [[o� -�    [[[[[[[   [[[�"\\\\\\\\\\\\\\\\\\\\\           ����ooooo\           � �� 


 \           �-�������\\\\\\\\\    \\\\\\\\\�I[[[[[[[[ ˳� [  ˵��[  �---[  ����[[     [[     [[   ��[[   ��[    ��[    ��[      [[     [[     [[     [[[   [[�pppp   pppppp          pp          pp �����    pp-----�    ppo-�     p
  
-�     p   -����� po  ------pp
  ��   opp   ��   oppppppppppppp�"	[[[[[[[[[[ �-���[  �-��̘[  �-���[  �-��̙[[[[[[  [[[ ɳ���[[ ɵ���[[ �-----[  ������                   [[[[[[[[[�>[[[[[[[[[  г��[[  е� [   �---[   ����         [   ����[   �---[   �ʳ�[     ��[[[[[[[[�F[\   \[      [      [����� [----� [����� [      [[[[[[[[�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                � 
               Y Y n r  W A T E R   S N A C K S  F L U I D   M O T I O N 	 I C E   T O U G H  L I Q U I D   I L L U S I O N S 	 S A I L   A W A Y    C A P T A I N   G R E E D ' S       