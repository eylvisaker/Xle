���  .b$
  :#>                          	
       ��d�ccU2�� DJ                    ���                  mq                    97;7<8;:   3;74   �������Q��� C/4                   ����                 kj                    D2��0//1K  H/11L  �������,V�� 520K                  ���                                       H�c�222>   G02/4: �������,T6   H24                  ����                                     93�ec�200;<L G/0/21L�������-UL   52I                  ���                                     F/2�f�110100;70/12/2L������-S04   90K                   �                                      D/�f�0121222/0///10N �����.�T2J7L9D2J                                                          C�뉏/1>@?//1/����20Lʘ�~-.,T00/2/02I                                                          �����1I  F/001�fc�1I ��c���O01/121/M                                                          �������  E00/�fcd�1N jutv������0��/A6                                                kh        ������88:7/1�cfdc�014     �� D�����                                                  mt        ������0220/�fdf��0116     ��F1/���                                                              ����1221/�fdfc�B/16      �?@��                                                            �   ���0010�ccec�MsEN                                    #                     #             ���  ���201���oie��dn                                                          !S4              ��   5212//06  idedh                                    (                    "O2K                   ?@5>=AK   ujut                                                           ?@                                                                                                                                                                                                                                    