�y+N   x   
                                                   h �`�0(
0h0�0�0(`j��`� *
0j`�`�*@l�����,
�l����P,@n�����.
 n����P.@p�����0
�p����0@r�����2
�r�����2@t��`�04
`t`�`��4Pv��p�p6
pvp�p��6@x�� �`8
`x0�`��8Pz�����:
�z���� :@|���� <
�| ���P<@~�����>
�~����>@�0�� 	�@
����� P@@�@�@	B
�� B@� �P	pD
p�p�ppD�                ����������������      �     � � ����DDDD��������������������������������������      ��    ����      ��    ����             ������DD����������DDDJ����������xDDJ�����       �      �����������������������������������J�J�J�J���������J3JDJDJ ��
�� j j j j � � � �ff      ��      ff       	       f       �      ` ` ` ` � � � � `       �       � � � � � � � � ���� ���������������?�?�?�����������������<<��?����� ������������������<?�����������?�������0����?������?�<DDD���������DDDD������      ��    �����F�J�J�J��������` ` ` ` � � � �  f j j j � � � �                                                                                                                                                                                                                                                                                                                                                                                                                                              