��N@   x   
 0                      P �                         h�����(
�h�����(�j��`�`*
`j`�`�`*�l��@�`,
Pl`�`��,�n��`�`.
`n`�`��.�p��`�00
`p@�`��0�r��`�`2
`r`�`�`2�t��`�`4
pt`�`�`4�v��p��6
0v����`6�x�����8
@x�� �`8�z�����:
Pz���@:�|���� <
`|�� �`<�~����>
p~��0�0>����� 	 @
����@ P@����`	`B
@�`�``B�� �	D
��D                 DDDD��DD"DHDHDDDD.DDDDDD�DDDDDDDDDDDHHDHH�".�D�����H""""""�.DD�D�D�D!"!!DKK�KD�D..�.��K�H�H��.��.쎸H������ff&affaK��D��K�..".��KHK����..����D�������������������������D��""!""����K�K�����..!HD����H�."��.����������n���&f�������D��fbbf������D������D������"""""""DD�D����""!""D�D�DDD����������ff�f�������a"n�����DD���+"+������H�DD�D��"����D����..�!!K�D�D�DD���������������!�����K�HD��.����H�D���.�������������f��"�D������������DKDKDDDD.�D����HD�!��.!DDD�K�D���!DDH�D�H�!"!"!DDDDDD��;;DDDD�DDD�DDDD��������ZTZTZ]]���������ZTZTZTZT��������]�Z]ZTZT������������DDDD����߯O�O������O�O�O�O�����O�O�߯��������D�DDDDDD