��N�   x   
 0                                                  h�����(
�h�����(�j�����*
�j�����*�l�����,
�l�����,�n�����.
�n�����.�p�����0
�p�����0�r�����2
�rp����2�t�����4
�t�����4�v�����6
�v�����6�x�����8
�x0����8�z�����:
�z@����:�|�����<
�|P����<�~�����>
�~�����>����� 	�@
����� �@�����	�B
������B�����	�D
������D�                  ����  ����    ����  �?���?    ����  ��     ��UU  UU    �
�  6j   
*�� 

"* 

 (����  �`� �    DDDDDD  DDD  DDDDDD