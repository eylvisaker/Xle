��N  r   
                      ` �                         h0�P�P(
PhP�P�P(Pj0� �p*
pjp�p�p*l@� � ,
0l0�0�@,Pn�����.
Pn0����.�p�����0
@p@���0�r 2
Pr ����2�� �p4
`t����4�v�����6
�v ����6�x 8
�x�� ��8�����:
�z�����:�|�����<
p|p�p�`<�~����`>
`~`�`�`>����� 	P@
P�P�� �@�����	pB
`�`���B�����	�D
 � ���D��� t0�P�@z                 ���H��ߙ  ������DD������������DTTDD���..�����������������wwwwwwww�������ݪ�j�j���������j�               DDDDDDDDUDUUUUEUEQEQT����������������DD�D�U�������#DDDDD���..�DDDTDDDDT�E�D�������D�D�D����.�n�wtwww�����wwww����tD DD�����������������>/^//E_|�T�UOU>/>/>/>/<�<�<�<�?�?�?�?�?�?�?�?�""""""""������  "
"(����#�?�""""""""������     �D�DD   ff������������������������������������������wtwwwwww��������wtwDuDED����*�B�t(wB
�Ш�
�Ъ�B�t*wB
�Ъ�
��  � � � � � � � ���y��ߙ�����������������������������������������������������������    ����  ��"""�D�D�DED���������������������ЪЪ��ЪЪ�D�D�D�D���� ������� o�����     ���   




DDDD�D�����DDDD����������DDK�����������DD����K������ffUUUUUU��UUUUUUffUUUU����UUfdUTTT��TUU      ��    ����      ��    ����                "�"�"�"���������������������� �����������������Z�Z�T�TU[�Z�EZUQ���������(��DD����������꺪�� �
�
 ��  
�����     0 �          �     0    0 0  �      0 � � �     � �      �   �      
�
 ��  
�����         �   �    0     �  � �      0 0       � � 0   � �   �         �  
�
 �� 
�����   0   �           �  �   0     0 0  �     �     � �   0 � �     �