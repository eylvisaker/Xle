�Y�  ��������������������������������������������������������������������������������������nkm������pkl����nikm��\\\\\[[[[[�c����������������dnjikjm��\\\\\[[[[[ ��c��������������da jkkjkk��\\\\\[[[[[ ���c������������daa pjkkjl ��\\\\\[[[[[(�����c����������daaa pikl ��\\\\\[[[[[ +�����daaaaaaaaaabaaa  ��\\\\\[[[[[ +����daaaaaaaaaaaabaa ��\\\\\[[[[[ +���daaaaaaaaaaaaaaba ��\\\\\[[[[[(��daaaaaaaaaaYZ aaab <=��\\\\\[[[[[ ��     (   (        eeeeeeff;:ff��\\\\\[[<=[ ��+++eeeeeefff  f ��      ;:  ��,eeeeeeffffff ��  ��+!eeeeeeffffff ������������+!eeeeeeffffff ��njm+!eeeeeeffffff ��nkijm++eeeeeeffffff ��pjkklnjmeeeeeeffffff ��pkl �5��������2nkijmeeeeeeffffff �� ����5������2�(+pjkkleeeeeeffffff �������5����2�� +pkl eeeeeeffffff ������5��2��� +             ���njm����52���� +���������������������nkijm++����������(+���pjkkl+!���������� ���pkl +!���������� ��� +!���������� ���+���������� ����nikm���������� ����njikjm����2N���� ����jkkjkk���2��N��� ����pjkkjl ��2����N�� ����pikl �2����<=N� ���� 2�����;: N ���          ���  ����������������������������������������������������������������������������������%%�@D9-	1����������������������%%�		����������������������	 2| >)�4�
�����������O��     ��O����  ��O��4�  ��O��4�   �O��4�   �O��4�   �O� 4�  ��OOOO4�  ������������*�������������������� � 4�   �4 OOO �����4�   �4��  ��� ��4�   �4����ɨ��� 4�   �4444� ��� ����   ������ ��                ��������   ���������?�������������     ��   ��  ��˵���˥   �4444444�   �������˥           ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��������������*
HHHHHHHHHHH   ۳�� HH>11۵��  H���� ��  H>11����  H���� �� H ����    H         H ������� HH�գ � � HH��      HH�� � �  HH        HH  � � � HH        HHHHHHH��HH� [ ��-�  [[[[[[[[[[[[   [[[[[[[[[[[�<[       [  [       [  																		[       [  [       [  �4[[[[[[[[[[[   [[[[[[[[[[[[              [ �������[               [ �[               [ �oooooo[               [ �





[[ �������������[ �����[[ �------------[ �oooooo[[ ���ϳ����������� 
  
 [[     ��         �������[[[[[[[[[[[[[[[[[[[[[[[[[[�\\\\\\   \\\\\\\\    \\\\\                       f\                       e\  ��������   ��������  \\  �------� ---------�  \\  �-ȳ���  -ooooooo-�  \\  �-ȵ���� -o�

�

-�   \  �-���o- ��ɳ��-�      �-ooooooo-�  ɵ��-�      �--------- �------�  \   ���������  ��������  \\                       \\\\\\\\\\\\\\\\\\\\\\\\\\�[[[[[[[[[[  [[�����������[[��������� �[[ � � � �� � [        ��� [� � � � ��� [         ��[[[[[[[[[[[[[[�A      
   
        x } ` d  E R N ' S   F A I R L Y   D E C E N T   G R O C E R Y  G E N E R A L   W E A P O N S  R E F U R B I S H E D   A R M O R      B A R B E R ' S   B L O O D L E T T I N G      P R A I R I E   S C H O O L   