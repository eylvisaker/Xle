��N`  t   
                      @ � �                       h � (
 h �� ( j � � *
 j ����* lp�p�p,
pl���� , � � .
 n ��� . p � ��0
�p ��� 0�rP�`�P2
�r�����2`tp� �04
�t���P4pv`� �P6
�v��@�06�x0�@�@8
�x�����8�z ����:
�z ���@:0| � � <
 | ��� < � � >
 ~ ��� > ���� 	�@
����   @ � � 	 B
 � �� B � 	 D
 � ��D �`np~���                ZPZPZPZP�����������PZPZP  ������DDDD@ ���������DDDD���D�DDDD�D D@D@� �     @    �𙙙�    ffUU  ������    ffUU   �	�	�    fU        @        _____DOP���������  UU          P _P____� ������    P _P    � ��________��������__C@ O�A�  ________��������              DDDD         @ @ @ @ @ @ @ @ P  P              P  P       �  UU                QP��
�P�
j  � ���������  �� ��@ @ P @P@ @ E @    UU           * SPJPZ  ���DDDDDDDD  @ D D      D@DDDDDDPZP�`Z`Z�ᬡ���
jjP Dʦ�E `
j�
�EU� ��P DDZ ����UU 
��  DD���� TDD���UDD@_____ZRj�������____�_����������       PP         ____    ����   _   ��� _____ �������     _     ���           PP @ @ P _P@ @ � ��DDD���������  DDLD� ����� DDD�Ͽ(�O���  ( �@�@� � Ё * ��� 0�0��. .    �� 
� (rr  �� � �( ����� � =�� * ��� 0�0��7 7    �� 
� (��  Bt B �( ����� � >�� * ��� 0g0��     w@ 
� (��  �| � �( ����� � 6p� * �tt ���? ?    �� 
� (��  �� � �