��N  v   
                        @                         h � � (
 h � � ( j � � *
 j � � * l � � ,
@l ���, n � .
Pn0� ��.�p � 0
 p � ��0�r � �2
pr��P�`2pt ����4
0tP���04 v ����6
@v`���@6x ��� 8
�x�����8 z ���0:
 z@�`��:�| � � <
 |P�p��<�~ � � >
 ~ ����>����� 	�@
����� �@��`�`	`B
`�`�``B`�`�`	`D
`�`�``D`����                ���"�����3��� ����������0��
*误�������>���� ������������  �     0    1 D�@������ @ @  @  ��?���d�Ofddf��� �d�����	 �F��D����13 "*�DDDD� �� " �� D&@f`f �����	D@DDD   � � 3 3 30 D D          @ @        D DDD      @ @     @DDD`Bf���DDDDD@` �@ @D@D@  `f``&f��	�	���f`f`ffff	������	&`&f``f��	���`fff`df 	�	���  DD D                @  @f`b`dd&@������  `fff`f	����	�` ff`` 		�������`@�			 	 	 ������� Df$&`ff`fdfdf�����	�  	 ��  & B&	��	� ��&ff D`����� � f`f f   �@DL�DD�11  @ @ D                        � ��	�` f`fff��	��		�f``ffff��	�	� �&dff  ��*				��� f`ff �   �         ���
���� � �"�� ��.쪨��  *   *�  �  W W W  � � � �           u �W � ��� � ��
�����  ��                  �������������    ZPZPZPUP����  






ZPPP U�PP   ���� 33333   ��  ��                    ��� ��                     ��   ?�   � �     � 