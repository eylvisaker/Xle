�Y�  �~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~��																											U��																											0000////																											U0000//// 			38888888888888888887				~~~~~~~33333333333++0000//// nim			83888888888888888874 			U33333333333 +!0000//// kji			88388888888888888744 			33333333333 +!0000//// pjl 			88838888888888887444 			nim3333DDDDDDD +!0000////  			88883<=888888<=74444 			kji3333DDDDDDD +0000//// njk			88887;: 44444;: 4444 			pjl 3333DDDYZDD 0000//// iji			888744  444444  9444 			 U3333DDD     0000//// pil 			88744444444444444944 			3333DDD          			87444444444444444494 			U(   (  			74444444444444444449 			~~~~~~~,++				      (    �(       			U										)****)											U@@@AAA																							@@@AAA 	������																U@@@AAA 	�>>>>�																~~~~~}@@@@@AAAAA	�>��>�				@@@@@AAAAA 	�>>>>�				@@@@@AAAAA 	������				\\\\\\@@@@@AAAAA 																												}+,+\\\\\\ @@@@@AAYZA 																												U""",\\\\\\ (   (     																												\\\\\\\\\\\\\\ +,+  			c���������YZ��������d				U\\\\\\\\\\\\\\ ,,+			�c�����������������da 			\\\\\\\\\\\\YZ """			��c���������������daa 			[[[[[[[[[[[[[[ -----------------nim			���c�������������daaa()		[[[[[[[[[[[[[[ ----------------- kji			<=��c�����������daaaa *U[[[[[[[[[[[[[[ ----------------- pjl 			;:��daaaaaaaaaaabaaaa *        [[[[[[ -----------------  			���daaaaaaaaaaaaabaaa *      ................. 			��daaaaaaaaaaaaaaabaa(*~~~~~~~~~................. 			�daaaaaaaaaaaaaaaaaba U................. 			daaaaaaaaaaaaYZaaaaab nimnim............<=... 				                     	kjinjikm           ;:    																	

							pjl Ukkjil  																										 ppjl 																										U  ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~KN#LNN�J1J��7IG�����&��  ���� � +�8'b<�Bb��������������������� �4 OOOO  �   ���ש� �4�    �   ���ש���4����   �   ���ש���4�      ���������� �4�      �   ��  �� ���  ������  ��  ��           �      ��           �      ���������    ���������HHHHHHHHHH��HHHHHHHHHH �OO      H   ��  HH �OO      H �ϵ���HH �OO   HHHH �44444H� �           ������ � �                  H �OO   HHHH        H �OO      H       HH �OO      H       HHHHHHHHHHHHHH��HHHHHH�(������������         ��    ����Ш�    �O��Ш�    �O��Ш�     ������(
�     ���   ���9/////////� 4OOO// �4��/  �4���/  �4���/  �4���// ���  //      /////////�#���   ���O     �O�    ����  � ����  � ���������+���������  ����  ��    �     �����˦�4��˥�4��˥�4��˥�������5[[[[[[   [[[[[[[[[��O4[   [����  [[���O[   [Գ����[[  ��[   [Ե����[[    [   [������[[���            [[4O�            [[[[[[[[[[[[[��[[[�A�������ʳ�ʥ�ʵ�ʥ�?
���44�ʥ���  ���   ��        ��        ���   �������ը�����������ը����   ����������������������������������͗����������������� �� ������4�������� ������4������͘� ������4������͘��������4��������������������͘����������͗��� ��������������������.����������������������������Ҥ� � ��OOOOO   OOOOO��             ��OOOOO        �     O        �     O        �     OOOOOOO  �              ��       �����Ϥ�       �44444��       �4��  ��       �4��  �����������������A                x � n d  S O U P   K I T C H E N  T H E   W E A P O N S   C L U B  P O O R   M A N ' S   A R M O R    E A R L ' S   U S E D   B O A T S    P E D R O ' S  T H E   C L O U D Y   C R Y S T A L    T H E   L U C K Y   W I N N E R 