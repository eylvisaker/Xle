���$����000�	0                                                                                                      F @ �� �     @     r��                                                                                                                                                                                                                                                                                                                                   �$$�                                                                                         �  �   �  ?�  �� ������ ��  �  �  ?<  <<  �?  �?     �������������  ��  ?�  �  �  ?�  ��� ��  ��  ��  ?�  ?���     �  �   �  ?�  �� ������ ��� �  �  ?<  <<  �  �      �������������  ��  ?�  �  �  �  ?�� ��  ��  ��  ?� �����     �  �   �  ?�  �� ������ ��  �  �  ?<  <<  �?  �?     �������������  ��  ?�  �  �  ?�  ��� ��  ��  ��  ?�  ?���     �  �   �  ?�  �� ��������  �  ?�  <�  <<  �?   ?     �������������  ��  ?�  �  �  ?�  �� ��  ��  ��  ?� ?����      �   �   �  �  ?�  ?�  ?�� ?�� �  �  ?<  ?  <  ��    ����������������  ��  ?�  �  �� ?�� ��  ��  ?� �?� ���?      �   �   �  �  ?�  ��  ��  ��  ��  �  ?<  �< �0  �<     ����������������  ��  ?�  ?�  ?�  ��  ��  ��  ���� ��?��      �   �   �  �  ?�  ?�  ?�  �  �   �  �  �  �   �     �������������� ��  ?�  ?�  ?�� ������ ��� ?�� ������ ����      �   �   �  �  �� ��������<�  ?  � <� < � <      �������������  ��  ?�  �  �   �  ��� ?�� � �� �� �����              �  ?�  �� �� ��  �  ?�  <�  ��  �< �?     ������?���?��������  ��  ��  ��  �� �� ��  ��  �� �� ?�?��              �  ?�  ��  ��  ��  �  ?�  <�  <?  � <     ������?���?��������  ��  ?�  ?�  ?�  ?�  ��  ��  ?���� �?����              ?�  ��  ��  ��  ?�  �  ?   ��  ?�  �  ?      ������?���?����� ��  ��  ��  �� ����� ?�� �� ����� ?�����              �  �� ������<?�� ?�� �� �� �<  <   <     ������?���?�����  ��  ?�  �     �  � � �� ��? ��� �����     �  ?�  ��  �� �� �� �� �� �� ?��  � ���?ÿ���     ��?����� �� �� �� �� �� �� �� �  �    0      �  �  �     �  �  ?�  ��  �� �� �� �� �� ?��  � ���?ÿ���     ��?�������� �� �� �� �� �� �� �  �    0      �  �  �     �  �  ?�  ��  �� �� �� �� ?�� ?��  � ���?ÿ���     ��?�������� �� �� �� �� �� �� �  �    0      �  �  �     �  �  �  �  �� �� �� �� �� �� � ��?��� ���    ��?������ ��� ?�� ?�� �� �� �� �� ��  �   0     �  �  ?     �  �  �  �  �  �� �� �� �� �� � ��?��� ���    ��?��������� ��� ?�� ?�� �� �� �� ��  �   0     �  �  ?     �  �  �  �  �  �� �� �� �� �� � ��?��� ���    ��?��������� ��� ?�� ?�� �� �� ��  ��  �   0     �  �  ?     � � ?�� ?��  ��  �  �  �  �  �  � ���?ÿ���     ��?����� �  �  �� �� ��������������  0      �  �  �     �  ?� <�� ?�� À  �  �  �  �  �  � ���?ÿ���     ��?����� �  �  �� ��0��������������  0      �  �  �     �  �� �� ?�� <�  �  �  �  �  �  � ���?ÿ���     ��?�� �� �� �  �  �����������������  0      �  �  �Z\^`bdfhjlnprtvxz|~���������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLZ\^`bdfhjlnprtvxz|~���������������������������������������������������� 					
		


 
"
$
&
(
*
,
.
0
2
4
6
8
:
<
>
@
B
D
F
H
J
L
Z\^`bdfhjlnprtvxz|~���������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLZ\^`bdfhjlnprtvxz|~���������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLZ\^`bdfhjlnprtvxz|~�������                                                                                                                                                                                                                                                               